`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
eaJ3jzLVN4iYHshjFGfH7iDwby1qtsbUgn9NsTJfPorjD6w/GWCOxand9k8gYdYsE8H8higTQQij
Ks8gerxQgQ==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VSe3tKso7/K8cXXjgmLUDRvH28kQKWXJ8tTQfX0r32/UZOwlNmxIePfSYtIWfuxt6ZOenjrqts9F
qDm1/aGT5K7d5lAisRNv+5ywzxaT1O1FljvvlCLsnGXhGOS1XFnkp+gyNCB8vFStTrgJQpWe5b3Z
eoX1P7QPsAD+pPu/HIo=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
C44Dv1dsP4amcta/a/2+OMbz0yoNp9xSsirtTnZBJ9ko038F6nYqqBn3ks/nNnutL+qyhNCMjsj6
HryQHGHqDTBPcTU7megvVzWcOpUf9VVtcG+ICnisuRIUcamMq6rWv7Pgs14O3arFIlYbDLZ7pGqT
rC+/E+kLL6eLBIxNBq5vJPFS0AZUUuy8ETwyjI+HwSHUXjC2+qCvodV3HgBelmKBGOFYdSvo1SQE
vCC0pK0JB6pLsdm0BIpYYFtBCK098p7RhkcsXgUTv8Cl5KkLc5J/yClw84CG6aujKxU6YlaqDUkm
WjZDlfMDf4YiD/B9vDKWzN9j7aWckcDAzKy0aw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fPe5Qn/Lva+KXqMIjztyKFNigW2k6dlpH/yRpbs1Yt3JMqvphI1MkrlEYtmNM05iK+bwpYz7K+yM
epVPFv8dS+JNSOILozSr7Q5d7zuzvVz+RH5KD5toQ7ZFL+tqv9biIsLC7hxclKccUUq2lF8TOnn/
Stfkytgww0uOxbNmLRNqb1LVZvqq5Yia/dsfHC1RWoBGdX/5p1PnNcv0amn+2ctXb3sWEOmL36qh
fcB7qdP+XVJiaRWXInKS2+FH73TIwvW5GMC8iqI4aW94fhoyt1ReENmRo4eIwsdHZjb4b3uPKNM+
ydPDscCK+XQB22zQWqUcXkPmfm1y7pX2Gexk1Q==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tCxzQ9cYgTsMBnU74brLcwgE7ZbxsKnDQV5ckyHI1zahUjRSatJmRev3DiXaUvddc7dmFgbdsIOS
j7fYTw4tqrhOIJBvQDePYBu3rc1v3K5B8LW7qI1ZKgQeede/k2r+syqrvQQeQg0a4fwB2c5mHEbl
NRZ69UrpB/PFUv29Hg5nYfIK7V+ODpQGXjB853+067Cr8fvaQRvNpAEidb8w7ye8Y6xHJBhxtUCW
IrS6xgq0SBTS3x4IltuhiNblTV+pIbDim59znmg9TY5qrde9W4juI6INcUfTXoqHFHuUY/uhQGqt
rHIjCX3N7TapP30u2za8+rEhXGGeBQw94uhOnA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o1m7Xa/RBgISQWxhUvD5Ea59hySkU+QK3550vwS+kkjyCgo7Ar3o7RJ5AM3ZDARWop20KPTRKmxq
Mm54cgZ4LvP2eVH94Np5QpRH4FDpALUXqWx+ItSxNIFep2ERwfwxPhcNdoSFcHaS3j8ySwqYLIc8
fWEoImUI559znJFkh58=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JXv7XsNy9y7hoWdO4Yyzh8PS5yfrshxXy/hSvzb3WQPdcLXhJUiUdr4SiUCE6m27wHxvPwTS2wYX
mEEpN+lrAABNfKHa6mVrMN5D2K/KHob/ENdS7zhbhMdGmyqPT4fi7c19ASRRv5hdRQ0gGdfEvH7c
CkZCUcUlurmoqVvf6jc/VOmV0TfpUAiK3lxnv6wNwT1exD437GwKQxEO8FJ9EsfkuoUilwl3r9wM
I/u+l7Rnwl8/tnm0V4kp5ptShgrUloy0f8cZg1r1yZ6zrHPooaHqWw7dGO4hwWmPl9756dNUXiIf
eldb4yGx8O1ES2HBB3sT9dByfFD5DdLtmqkJBw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 610096)
`protect data_block
kl8rkJWDSsWNTEwjL8bz7I3usy8xlDMv7JgKMo9+VwFoPeGGZMdMauvj+F3NUFYHeBHWGviYrBUb
Hdism9AgSgGg0MrGsQAmEcDp7g0tJVNVolOp7EQe0AVWd3v3xu5osn6/u7xs2KyJs/m4t1eMmcP5
rim/CAZRgY4AXmOG7iA+cPMc9vXOw2HNqebYGSGN7Zu0P0Oa2ozG7E49IcAt3BnGoP+Zy0itJ2tu
gaUzynx+fzIGIm2hppv5aJu4Kc0/1ZBAWAmH/QXUTNN2VRt3VVSa2wBnXT9lEB9yGk3jMbm7ssrS
45OPJx6kGD9ULe7qafgqgrh9rMcv62T3T6aCyA669D1ntTZ5ssnk0Z6QfmmG6VfHFYeQq5WSrS5V
IakMCG6dMgtnfYgftjC/+EvzAYBuyrT/1jLlChc3WmhHNUswVKaYUV5CDupdAtQjrBS8lRxxRPT5
QAIcfYYG/Fxzqn9VAyCMNYxY70wKYkp2QCdBI3o7HOQJOzh9dxpfQnPLq+1Pv5DOp95ubkZg6yHJ
KWNCe+7TORBhaI/kdsOHIv4loSuwvr30WliylqJYG3fowqSmMVoUxZQuwnqEsPz+6hDYcCtdHJPk
/TzsyAEXi+irWy4E+uOsPsj3uaKtu349Vg5dcxNIG0/MNGsunaZ4+/YJTXNc1Ux9n+DTfcrP/Bto
thVc5kuNyxlzEn8hmgIw7p43L1UFql0hRJi1crEZFA9TJeEvaZvplLaFyg3WlqTY/0kO7gNyMEvG
6J3iq/XhprK/BlFmYbUXafWHC9a61SujQCWiN2jZsUsn/VEWTQHc2eb1o3VCzpdzPmAWmaxvKxh5
+GYg/1TMQ+h4k3RKCfK22DGJCA1VA7G1A0QkwAdlflNajvv703xHRyHeU4sZk2n06YNK0TaLy67z
7A+9Wo7N9wYr3ggoKGDoSv0METk16mnibQBut+7SMkFkqOZ4nTldnIwjNg7YR2NEgVdAxzdxdAMG
+wLZ9G+2Z/ybxYnR+IuGiZ8e8kFJetpS2ilh2Q4wM/LbcpqZ0pIjTeJCr0es90PJxe4FlIJcv/b6
r6PPvYXjcxYia1T4sqexlBY/tZqaua+wfjUqoPziJTju97PJYI8c5p5o7rUf/uqhtT3iDcgGcGhs
xfGmLCiJ0xwWuSrOX6j0HHq+VdJ6mOmS5YsbXTmBiOT9EJaEpdNYtO9+tB3CCVOVXPcD0rXol44O
fYrooFldtbyTOFIBOCUKrBC6Oe7efMeSHCaXt8QilS7QvCN3OLXh3bTaH715IaMlMziuLMA3ujIp
EXsdTkFEQKJ8OlHAQ0qIpyAb9t1HKj93122EnWaFuIcVFNtL+PjihczBvSWiLkwg61NJkhc4kBDg
GUGtA0efTuvCgjKW8375zAZd55qyvVKzqwOQToEsJR8gK04oNf9fJYYDvC+hjiINyYeBp9U1lM9L
o0QD7qkcOuOF1d6OhPd7umt836hQ/h+CmZ9/BwPdRFLClPYRk7jhzFjpEoAYafiJWvH3ayZHCwzD
dCazRkbpFmPBx6Ur/LLd1N1KAw/QE2RRvl+BrOvEcsHKCS2M1TCruH+H+cud5cXwS8rgrMxR09ud
EoK15sIsXizt811TfYwfGi4hTlZhfuj+MU5eA6p4UgaIJsC6v5Vf15gXMm/jHsUEy6dQeAtxVg1n
L0knTIK3hsCYIIXQ6qDw5EhDNHGZEY7v+8r5DokMfWS3QVjQykpkKYR4oTn1jSGNFC9gpUZeX8Oy
owQ9x3Kgu4/ohdXDWxsMHS/Tw6uElAfx1joepBSYmuf91eWnExL7vd4NalILJFx5nPpugwequE9J
Ozf/S5YwxdVBoWEamFDdQFXlfRVdwda20BJaxw3UJZfsd/eGXiszPsQUGNK98tbe56kbY6CQZqFx
6rwKsXczqbp7S/4J/7QFKM5pYHY7NA27DcyvsHygNIK/huNn4a0Rzw2ZFxJGxHjy8C/KZKRSaTOZ
7XUQF/LXh/Im/YYJU0kMWUAsVJRVZyAfcsPJlVkfxaPlCXYKJJ6UP4EhEjYp+iFXiqZP9w5pyMKu
xtPneKga79KxeDhEVZQulnvkRCxNPkd3p+qGN018JEXSQcdQb5MK52Qpvq6tlykJFNHmBDLD59Zc
SXcWk02GSnf2w6NJQVuFzbD1G+cHAPu8DG3DcB7BJDrh+W/Q+pDYySdV9Kv+u3cEZu3U8e8HKV8H
CWi/nYR4dUoHFP1wxB53aFDvFnMBYKgCybnxtck2Ms2cZTD2NxGo6NhKB57+MU3GM6KdSPxynOjz
IG03fn5tAb9g5/1+H7Naq1kFj6mOLKeJTaRi+GHWNvDqibg4ASI3/9PehS9WKr1P46RJ+YbSWDDD
5ENnYjZJQ/YhIrE9PclslUEfheelaM6K3UxXomG7czGfipCERNt1fgC9mCj68JvDYU6jHNrTz3qK
314ZYSeONi0Oeje9fkKIAMXABxiAtZj3hOOVHEECt4oQ1Ri7SEuu1IfeqHnCfkYkTL6fTHIqbmuM
rrLp26UYevWhp0ptnuIqWq22oP9tKKQvq0k/kjFrF/B0iKoVGVns92NLnSjl1xulyf48YevX07ZI
YT6jq4wy+fy1ADiUE4UXMfgY+vYN/F3ULUrYjEpZ7VUq73NWi92yIvcVu1UUfyw382U0FFObJDRN
FrTMjKwr7XTtOrQTP5m2MT3oQUAz+Mxn7aebTBkBw//FzRlVTvQ9Uw5Ut4XOU33e/U8vxnE/Zlsb
lZCVEROCRT95oveSQz/BAXdevldxpJLflQDjfMO42fBZRNzc6hnMemPz0CgL/0u2R+KqNju+lNNo
24UhJseP3v8EHiY3Ho+kRatiofoORaWPelB0xjFPEQE/u39zeSydI2hwa/Udi9pSQqjxaIspwxli
mmQeygNzDr0RWUrrvWUMcDgyJURVlycQzIriDAOD/rcCGUI7b+2/YZq2phSnUmd6Gp1QrwQX3hjd
Ad5UQtniN8/MqOswPqx5g3+vSjJuaZ7vQNHyJgxstbOCeQXmyN1LN+GL8y10d7y9q0xadVtW1ksO
AT5uXQj0OeHBo0bh9tVHdZ0ixpIzgV48pVFNWpa339EdQjJ1nKnYhIB6kYe1y3zBJ8F3y6f64BZ4
I5UdHNcvyPLgAmgn2iZznruQMi1nO4Xml6MJvsmAKMgSX1QcmrEWO103SPNMt6cgmjq/RrWvqkF4
ceOx2zoqYn7j2mCMtyq6twqPIF8VplOTAb9Q7K55ntL/4ggOd0UWfcPSX7Ksuj8pZk4B/KHKsqyw
SkFYmU3ENYoFw12yVvC+0mt1yaaNRjud5KDzOumSwhd0BVnxyz9q3K7GGyEm8yX2yYuIkiUznMhM
A7ac8NRvHGm0+K0xLghd4urjd4+//5Zh/f8KkTCdmbS0QOPzW/kFNeuSedh8jHLCMSGre/ppf/dL
jPA9KHQp53n1hKOI7WM+4YnERtbz6zFTLzVuAFOLVN3beFNRj3OHcQd9WsRdkn7+7B057Ayo4zjb
dkyf+FYh5rELfO2S7jk+0bAehUaDsoUNF9o5UUiNdiWJ3PNTipoVgGsGkVM+yJF7zmT8JO486tkv
908Xx6uCPbOTVATpJ85rPInV0xVRGLvuT7jQJM1zdHPlCHGTUC+5AmLzBlldsZCghaugfMkTUMHG
yYuIVPEh1tEXyCqdYzTH1CTXBYZtEeP/3bV5BO2FzYk1OXghTqsjDkO930aKY4NffO5iR/3TDbhL
uxWw/8GnoueY1loAlY/CCGYbYaargPH2mN44uM5cE83m/WyVYYFTSlw1PvZ0+DUpXY8RSHjP4uDm
3u8fY+3+UzdyXsAQmmaEo5dU1Ayy+6NEHXFnnz6GoThk9HdjgjiLKoE71trCB//ZzX1ujJY1yIsW
So9aQHu4b8HksLVaxyvwLDTnW4ex/ZdYgW32UA/DERLtRUJI2hGKSBZgQwkLSChw1usYOCmEVXbC
AtVV9yoDX1y1XwEe1DPN6iU8A06ZlfenQBjeHtWu2A8KE1bvhFJfWigfUUhJIDKjibcY5ur96suV
Y8dKQxj8WR2bdcJ0dadymvXyt05ifxXN0uBP+DO4oOypt9K14gPOCMAGvPbsQRGX0T316MAlu+PL
c4dj++RvCHo08l7qkjdoorS1ekFXhyLRNymxT5aKlws3DxFTanAetCZ4kEBO+/x2dLFRC1ISsyKc
HwO6BsMzZ5y0lKUFvcVdsDO3WYpX/2lUr/VA3hLeAp0+7ODe692GlPMiwlfA57N3Jdbpzg67qP3A
AQqn0O39soA8bJAiOxcibZZ3G3ZSthXKTGPZRSaGayrvGr+7vboKgOjFkTmsgOXQJnNEXJ75BdOz
0zTncjtoFy9ZZnPHlpEys74H2gIYDgPfM1ud2UzA0EzmbjYSVM75QQHKCmheHaER3MAvlI4SEfXN
qeBisHLkP51pNUKFdidpnCrmkAxjoS8AGyQfkmNSgUtlF1mOiHf2PBm4tPE3kavSrpUIbEQqdU0c
lsZGtqhqjxMC4++L2PWNo27+SKFYU9onynhuSN7mRtdSp1qCfGIGnWAo4TtKBbTV2uIqbpTdAvhR
SVMjvqn2a72sNk7Vx1fXudiiDhOqZVcO5L9SlQv+w0T36j4jj6Vk5w00D9u4UtxkTV5WKH6Nmwct
uvOt+zTA0AJjOi5wWdwNPKpZTf3R2oFmgYMDr8SDvB3dMtD7w7tTWJcwDfHzl9fU56y4/iWWrpJ/
rZrtW/AaKvi1mDe568CUrI1LhBKgraNLg9jjrJxHjJn/odCFcU43DWvfuu77VcJmAnCSK0qprgUL
Cbe+TFrHYvZ/2nqIgWOZubCDeFZSsviwiF5WFt9Ov9Jznya3PiLBJ8/GFdRsxacPrASk3kAivK54
nJpmA2EF6DNBDLIqJMgTM/XqQU1xXtz4cHHl8Cz3xMbEFowap9SxCTITnz2EAlaLtJyseTqcPB7O
TX08mZRRRoBjRYD980qjFNkZRVmkouaXQQ42lrxghflzfKz8CAjNP/9eVWDnlE6rHZ3qhzCiu7uu
5B26gxjHAfUirSf7po75I9Lh6TVM2fdQGs2JoQ45R5v0gDLh8mm1JCiz5tu8yW2EpTQvTm+fFE2g
Lc5ablP1z7Xqv+K2SWnZf1sDnfXvaeNqKsfMn2rQBzs45rjHbvujqLyYzrVKKU1haE1lDKkPfmKi
exRlu4kQkGfn3EiaiPws9gvG2IdnH3wW2rH3hsHXNnS6jzJZo+6bWXbHaDdGx1cbcJGHaE9cMV1e
LJAPOglnk+AxUqnGJ75jrz9UPhCEb/Sx8dGcrwghEXRpPP1sOabrD3n20k6BU6gfr0oNgDx8TDOH
4BOQ3jOaLntatlAU0WuOnytpZ+TGw9g4DuyanSoA6Dy/sC/k72sVxKQUb1S8cRlBu3hqJ56pizOL
fQcCgVl1e0egJLkRUL6Yn+6G1VsxbHQ0eq4gSVfI0ejqprwmsEgrF4o6xeo3Xj5rSzAsBYiLvGjb
aa6aVtiAsCUKQBdmksTKrq9/0HW5lr1gnF3A6zXUMcDZBxCiBfwwWv7V+E2/M+RSKpYDpu76Cbpd
0DHMVD9pphQdjosZiFipqUlZQqfVfXYt9qYU/35dTlMBimEu2DwaKu5TRNgtJ4i2CDULPWPP7VQw
e64fHyyCg1P8z7IVFnJ76l2yrt5i3wyp8LSAdQKZbd38ZbNeCUEzvJXRA3OgryLXb1z1JyEsihGL
gktvP4Co7dUgW7ZeNyU6NlX0soZ/yPqs7PraNfO1X9mNEpeYfdalEA1hx9vHQ3xfnlAiDiFm8h2N
1ULOadvv+x0NXNbdKzkNW2WP4ZEufDcRZ/dNSq/UbsOaSg80JTbcmdESTN88jAEPN5ycaQKy1ELb
dztLcowA+5+6v/0O2p8sahJNPsXoCrfaY57oIIRT/kkuRhQLSHfd9/T47uqlrU84faev2tuKMAqF
nX0G+HwhIieT665KwwjjFfEUFOL1iF3SkwHAuTX5M4a5PKmRZCzMIeFvf+TNMCw4NQdcLoZRmdTX
9i32RwMzZpzGbunotcStV58mCdwbOyr3xXK7I78rTrhKwvG4krKWfzAJG9UHkQiAPRJTFel5809g
ujPZlpBLy9oYTMBAmKLTpm26jxP0qk++fSSr3vdCeFPN+30VAU4BFmkCNRmJ1/OxT46MBMavylPp
jQPsgmmez5crwQEnFRZaE1mpcuJR+GAh6rW2t9C8EK1LfmsDe1Fbyp5YwOJpqbw4dx3Im2/TOeP8
RADPXu/A2DWG3JQf/N4Io8ZmnfBgDj90E+wge72ZPEU0LejDI5/+O1RIKIohSr+lJn7hIa2NmlIH
evs5wYcF9zfL0mnm8O9larBc5WmdIz7CSxevNLlo8bSE0G6kVQ98A9M8jEma/Fwq3cukUQXSl8FK
yXVomQHQScPT/uK6D4Tyd3aPbJ98hH6Tq+O9e985oKyNyx42lNJe8j6YZH4aRCa07VJ4opJV5Ofl
JBs05epvc4affVO6AN/hDIlX0flmcDVA2+UNwJzPADZLWFgQHHP4yUzFGpptMDPP8P4Jnl3kR3Jr
1WbpQ8/qSwXL18BS6705ZpCu7b3MhEf2yPuzajjc7XgXUQ40U/rMTsijsd1P1KD+hSqddSeQN+wy
6Z1Wqugs6gmas9X+qNHB0Ipc7GbmK2K7jukQpcH1kVXdGhXZdeST5zlg34pS5cCelxK9wLRJ52hF
+cq0ZS7k+6bQP3TrR8p8920genADhc5LcFIE2XjXYhrnlHuUJNHpuG98tK57Qfi26vwsxGcCwvNO
s3KIYg1hYDVJAna5NbiWOzbXDKbOVLOE3MMaViXUUO9w7s+BlEUeBGrlya+f8Sgb5Xbw3pYuPsU8
VTin+Cc9qoKpQPHSTrIK/rI7lUEiVJXCgLuleupIEDLxT1gFIHQQwsfxpbfXcPoh/Pbm+JPGQzLZ
r0oShaD3bG0Lv7YSyISzG1jsN0EiXF+f2ylRvfpcYpeIn1mmQuAW1mST7u137hxlT0QsP8tlLDJG
zdU/MAGxhKw6R6kEP8E7hp25BDoznx1w7JhTH1FnR1JpH+yPmOq7URYnEruz8n7KkT2qn+Rdgjg9
Oj/cl+IxrezRMAjme9fQnUlP8BrlIs9scREWXjxHZBX1zZ2njnwqBKC1n14E6W9S9CfItqO+hbgj
VIq9BiqIWvyXkOfXSbkO+hfd4MSh7Pk9o5lh2Bvw/SdPE41P6uJR3g3MBm3Sl7+WjIY6Fh+hhC3H
2jhan2gmwaFW4XUVJp+79CCrEKwkd3NWWj4ye0APqI9bXW0oTut9xxxu5EWo8kpFBPM3dNqrxyJt
3aFqS8mJBscAwyT/vh3Ou2Et//zBXWCLVQqukEjZFxYP8OUqdcoQuTOkw3757qGpBs9tJC3cqp40
LV6tuek8FmPSWDsC7HOJDRD/UV7eqNOvY0lRjs3vXO7NJgd1uyTlERkxFnQMCFa8loUjC46m8RZg
O3JEB9GvXKM4kg07RXG2JwLWg81aJ1iF9YsHuboVp7I4ez2l/83SyapKw4+cHUA9GlYY3CpcE1o8
FSrRkghf5G90UySL75flocipjsSdNSW7YI6PM0zVpfyA7KEZc0d35LF2Z3tteyQ/ESu97y820MLZ
bh+WbCkYgxRZOzd7zmTdrAeKFUTXd+AsP+KBJqYosQzc59GPODrGHSdc7ZA2/eeNjvFyWPwvcC1p
3Ts7BjE1fk9xNMmpLMda96E9qOKZ9mesWYmekSJww0N/btqAddhfL3GzQhBuemfhQ0f1pZ4uDMRj
WoRLQf9CxpjbeOE6+mnFaLgtw+u3L9gqdd/aOR5pnvw661eYWCaHGWfzM5RPDjYPj3l7SzwnKCC0
fuCm3upBHheKYQA0whbqM+xjyhyQIBU3F6CmGeP5v7AjGuG99fqlVOVirFr2Y8IPdohuiXrMfROC
qvZ6NRN+nyupBxNe9LueGzoPM9rvlVmtgfwUf4PGhKGHO0i0cEYA7dXtqyHbXz95hfP3q1KJT6QK
HynwaamaCkGN/F9bYqCpoEmRdJnjPw7bkaA2s5vEG1eSfBlbT85xHmHBxDFM3HJGPAiXSGchPrtM
npzAtyLwHWsEbBJlAcbt0Fr3OYXQbqnLXM/7evkll9e4pMoxwi010kOqsr5tVeZP9+N9XT2+mDOu
0+M4JJHt9QLA0eoQmSstYdLwF+ELKSM65DGR7iX6/AmJR7velcBoxZ4ylL/Xq9qPwxz1JtK2rGrr
k9PaAP85Kgk6bpT2QbnRwixguIm4qYgchSOgiaFs8PRZXymZNN2obbf+vyTUQid6FkyKhHz0Hm3b
L0fHvwJE6o672LAe/GoIwTsY9XGAaUrzM5rdKYteIrDlzz0tMRD3WBP+e/o3inhIo8XVlwFr0NHk
eY2Kvy7UmfIb6uw9tt/T0fX9o045sN9LKkzK1/EfrCyRBvYDrPTPhv82wqFJKFkTW26dNZQq6k/S
R5BLQOjzbvCd+JqNZoknhDGIZgtLz3JZcz9/co6USz4wCbtBbSd0qQg8i0RYxiBUDhL9oyIcgK+j
5eBNEQkCjql3xL4pgfo76OqE2mkLvvHvD6ENm73docv8xbpp22PICGmLcYNz64TEsvCm6fT8Ux0O
0x27QHo7TX13nCSvuVrXkY/lLG0uv+VsxgIFc8izUh/mFg6kJ6rBEu0IsK8HAbFusDl7/FFc/QYw
yRPPsugT8LHGMiDxclhL4LGbIV8t2L2WJ5VQESZDo/xw+y7/OTvdxA63LQcymdw+3TlbXDDiJv2T
9iNF+A3yu9rFLm0qomUxDpHB70HFPu2WjWPDIuwUCdT1KBx9eP4oSm7CWL/XAkI7j/tHxCUq1jRz
4+EV9XE14NOycuCygLV1dWq5OlH8U78NYx9IkX/eFn3OYsycNgGGwZ+UFMKeFcYCzEbt4VwrA8f8
HyRqLx5cfXjedrH7HSdeaQ3tEyEQaqSxB400/XxAoWRShcHzJ9hTgvssHBGf7c3l7ejw4Vci1p8i
0o6JTQqb0Rs78f0zMjSo0br2YxrugQjx0NCDC/nWofXd7QIIJYN5IAnW4ALOjqpCvQRx4YJX7y3u
mhSVDJw1LEaEENAzMP3xuM3+8NDnLU7eEBXxTaA6RDyyAC0vhJ7m6TACCqXbd6Lc7pK60S6EHih8
U6qUZXo1xzqpkmXwvvLkFLbr9mxCuapNF2xiCWYBu5zUx5g1Ds5ZrHlMe0aJ3nq63Wr3t3UVj1N3
YyhGtxQPb8ulWGdx+x4i3g0kiO/hYRW0p5nHV0Eil8OC3xEJoSzR7XKfDqOzpA36nR/UQ5NSYU/e
NB59ZU6vdysKL79oLx5UoY29HsZi8Z9jBMRrVEjVF4Oq5HQSSB6l7asbRHrdEHTAn7CMYuROkPil
GONaVMtpKPbh11tJZG9Qw4jW1FbkWc1g9k6UtSkjXN6+bIts0ReagRSEeKKsmyQtB8s8UGe/9MaD
70ihPzAYMXsfFFvN1CiyfF0cHuejrvdZMwYGxVadvllrATHyhwzl9l4J3hDZg92g9hnn917oDPSw
aATy3teC0zPJr22+O+YPJSUsGwBy/7FguUJP+KL9NZj8uCOs1ssXNCKSPAWigYLA+zcNgXeWsRSb
UrxfdYbEebQRGz8zlsAq0wrUXEaaJpZQLPnJXeHsTw+iqWmMK+/TKhCt7FW19n6Dzq2H5hBGXHOy
TdxEd2F4DcuSoceG+BRcrBMGIDWfWsW3uP8/XvYLz8Al6KxzytJM49d85qDiSX31PKZhijDtfoWW
z1uBmh5/mEPN6aDuSn4N7nL7SD25qSO2bGORiE29px41pcwDY0e4roXKCUTRQtkn6pjaBK5pf9zv
MQmalhgBIdQ63hOE+Zr8pz55xlyC9exqMXI5Tnn21OWQ3vepjiaMQA4kvw0ubXUWvGiyvuL8zDD6
ttO12OufP97Lzr9HvJdpDF+AhZao/EdtEPl7URBlowCbtS4rbGTL45y9NJ950D/GtbBr43ppBPzm
iOEds430e91+sWb1XWm8MpjBlzFLi8GtkPhI9grOmLlogl3f+BA6IjFsgTLWrqSgKhOMt+6r35qB
MF2DUjYtJNc7OH5nfkmD0QLcTQNGDrEhFgXIBkFRIfqOatNNMuCkjxqorgMxbfbX2J6DIrDRaFOS
7153TOAmWV/oy892jm1yQVXY+jinhji9NfKfj1phz9mh+j4ht5ZA0fzEMoIU0wQlBrQr76RypXeF
KystOX8h0IQrLyg86omuvgZ5ZJ9kvd6tZII+wVEYnthGMw4fuKaUUpJIcHqFowSR+K+39q1rfCM+
+l7SWf2XBuxifZ35gLeAFx3hhUbr45stDvazqbRC9s4eXOQTJ7zLJmH09+FUX/S1U25LICMQnKqQ
JYRl7/LcPpVpuOAShJWsg12zfz/x9YzFnw5VPqgnd3gkGkVdjz9rCYtUmMRzyVzDsDX5cBJe+IHn
qDw+IDJ6a03BIHN+43AFZxTz131R+XUskf28auIKsn22ji3AkSldfs2T2raqcxHLJC8/aYGjXhx6
QadUMJei7z+MTaibDOuvvVhtJTIfNe1LoQnpOSq19bnJ0vNQIROgiWa6XPVfr6w+bUJVRU14uJoK
fkwHzUbFv2Y/fF5cn2/3rQ4nK/8/hkRhtQ6mz3jfxYpfRByqDo5W4yUbgMwUx8bQO2Bv76kG4Adl
9n7Tqr5Nyc/sAd5gZmzLbeyggciiCq7mA9IHYtVGhlP+zEwFustxTpstOvvRcmVD+A+2+GeRzNlF
DjnSIT/2x4msJuEDqSSjeLmJIBnUlzEk1SUzDy8v+orzrJIhNeOZxzq05G4RUB5yH2EAZMKegZZH
ccUaqUX0bsucnyXpkOdCPUZPUOiTOVgLiBiFY66g1q5ny7nLDcco/r/J2p2lmmTDdvJZ8exnPbsU
duRnbhv+N49uRlxTCCX2Gqm6FeSoBQGBa8L+ADfh4xBmcEar8qBsL6VdTcBTd5QoNVpFivJ3ZiG6
d22n/+h7WUimqyXe5Hohtz+kW0FyJZBxNG0nQGKMTAn8M2oVcI+BInc7HmM8JwZMgZ5ugiX+ZCGc
bQG2v4KlgXQ7epHiap5btcRaCmjjaOtXthYU4J3AbOtnUh8aW52rk/yH1Ym09ClEfe7ICjsSwLYd
n/DxVr8AtR9b/HMgpCuhMB/L788YtAwvSahL1tgnKpD3/u0UFB8jRg2/rFynLWarbMv6DJAOBz33
JO1U1ouUhJ+0z2DlDMZA+doklI6WisWaDW5FqIPMCD4YMjJ9fvQ8XKxL5GgN3bLow1zG8ePRijtb
3EvtB/RednBWz+NMRX8/l0GVQuiH50U97hxdTKUrcJwq3ZfIu2NLs21yrG06MA/c2gvCgXNkvlZ4
l8RQoCUbt4XTO7Vf3e2KRurZ0x3UQkUS1qxzbYEvXwuTV/fvLiVu9WRlc+o22ECe56M57KjBwQYp
ka4edOnMWbihChKLuhA+pGqeSmrQYjAUXfR9Bp8BP2LrYXkim4wLURw6PuuBQG2wIIE69Vu0wD9n
kShhoiQGpg233J5SBKxa0ZI4radJHAObQzK8xCOUzFtjNwt5SksENOXQzo13cgT1oJ4zHbG7Ywd5
9SG0hJJid0kNJiXxhLTaqaFGZX3jjT8ShfNNvJC3cd7CM/YQJSwyglzemY/Qjn+pTPv4A+RNhVII
qp4YwQe3/rxcI10MROOtEuWmXImXET4YPk7JFXAhVELSy5EDsR08NmrTFuaEjBystihtRvWPnwRT
oIsoHrboMnNWzDyVmwZX5OPzr2iLv5wHn+tjnhX4+rzQ8oMfOmnyz/qttb18pDWIcpKdYLYYICMs
PLGS7yuDPwNR0Kq+UlWUfdDRRmc6WcGL2e0FjBeYL63p6IqK+pxHKO20JR1QMvU4O9+nhg/IUD4L
ph6Pd40RNt8zXU4QWiYL7yEQn2Km2Yn9Gumh/AYGLMqs8/yco0Mg2bdijxISmqIfRb5EiZsOhgT7
lrlvhWXhXWpnUxcQkRBwnBvdwrddA4tJhWm5rVP5E5SL/UcvdPuEmO4bGkEvFGrjfHbiMZmdfCZD
fQ6JqTtoebQQAE+gPyWFFL1kDhQQkS/zwWNTcLL2Gje4dpOtv4Xz/yABF+Du3JzaJviOJSYOXApm
+78sDe1OdQm08y6H0n9r9JDrRegEzrtCM9VQS/3BH7PHtcwUeddewq9Vz+kcqNSXvMivHdHlzJMO
WIuAyZ6ynKooBARAHJR+UkQ9lNhEZYo/8a4SceGMQIkPGSs7fkLNLZPK6+M36kZw6MICe2c4v6Ca
eiRTlGmxlw1l/tDztKtfNGd81yG1NLkWJuYLK++ixsgLbYs9vYMNZR/29+BVXlMh84m3QtiC00j1
zsUhtL/au7HokXn2drJxkfG+JxFH+oCYB5biIUi1mCiI+ugYc4Dh8J5V7ChtVbgK3Otk7KAFmnrY
jFu/14rxf0EYS3yJPcY41nx3q7Rm3eVKqfkrJFLre1FdbB9ne7aaxGvRxq6qeMiStOekpW3UhA/Y
yDwR5QkEsiOZ/iZuvUmkJBcygo2uYCMZjbSJpjn0MKZFx1G27XIBMvgItFCyubtwrC0aAE72OQSK
bZo/9Rbp8rCEGASHo1uJfaNb8NaytgONLceUHTFMWYhSMETBO6mnK1LR6MXNbWEJlBBoBd5fH3ff
JwD4Hmz9BInp+gqxX62KBv0Td1G7xpn8ms3htyKEKR75U5owqAyAcxBqPwP0HVAiJfgG0CZ4wfKU
Bzgl1ESIBNQ4NlJiBuitUIduE0j6P9UjpkkCzatedRoQrcOwLwNOfhbBhxwnXSSAPZTzQ1EulxBf
Ztv4FhvG8qQJXgogOgW/V6jzBKyMhirfExi7nwrcRTnFqqu/bNIt9CjpW+Q0IG71i7LXfBEdAX0g
Xd1C7H5DEXZdJap5eV0PxH9bZxoV1TJiZuiPpTr2gu5jPTPoczI9zcZoqeX2ssKENVncdLol6Qcr
qRUoLCq26gHtAURc79i4YZNIEIZR+juaKf+BpEtC3eXTgK23q5jXKq0IF2tUWN3Zz3hhi3TbQt2u
493JZPkwSmxCVg9C0KPa1S9/1gCWjd8qKB/IAVTNfkjChucpKJXQv3uR9c/v1BpOKWcSCeKwem1m
U2vMYRPjq9tgQeUelK8HDuRpXhiQAWgkJ1A+Kf93xxnHTWA0Hr+F4O6jnVg8UcJbybXU9DljtS3V
LT8fRlo9QU/ixNyOCSx5aj9VjctdCwCkpCdv/RPGtNvGATT9EjqOJwR0LY57QbddpOm2pSuQlBbK
tobCFNVAPki8k6BEtO+HMAlHX3jW02b2BWEjNkUpEBx4oB6OnsAlgWd7x6RiJO58wbx57a6vA8Ln
1F8vwl5ijspbcIqN7KKvsdF/mQ6A66dxfMfQjmpoMdZtjXWeNmFguwve8l9B0ut5gXuKWAEUT0ZH
nVX67bE1cKiTzlHxyr7B91h2IV4bc9yMWOwaQFD5cqnkKM+Tvr/nm+fxdM+xVZXkahapFk5UEuxS
dhoKeqcx2ELt76Dtsj/+clN1BfbIDkGktg51JDyA6LXHhRqmAlFurIIKGJLKEx/ma5zjiVf41TYp
0uJmCnCR1ci6qYu4eO6irOR7NukS7C22qOGujcFmq1VmqIHRPUPHMP1Y6MrV2S8GawpUQbhQl1ji
MY7FYqt8T70ujEd2v+nCqEBgWH805T+Ie5d5+H++jeNB3P7W+2xmx4HL7O/0SJZRAjF0gdycXBG9
TbZTixr22PoTKLuQrHJzECeCLBFUAyCm2VrUZoEWMgpthAGLH5u8xXcfhJPkrV+exvV5H/xkJIb/
e4XHlh3QmA4wH84ot0sA/Hec0iowp0Ex+RdFlnsdLIE3pVi6lbaLy6B6S7+0c7x+cW+kwADvaYf6
OHVbxDi62W1/yCBZrd/X5HXEG5NM7ZD+Z4nThKmk2FsRgL9UtAgG1UPij8XSwnK6kw+T6rORw8I+
+neEEQYwjEcsC7pjCwn3fOqxyLZIWawO/IPp+YZroaGrG1VIMcT4lrst4JUqD7YMQbg7VeFo2Kbd
oHzgxx7lpxryWLUS4lYR06TrP/J8YG4MvQ9X3dNtP0QEnlyQBKLbo1tIqxJdP/BeugzSuTZ6xA3f
v/ijccpBOHXo2Gi4IA8A77YJm5mDfMCODP1J281jIIvcYXKSjmk8Hoo3bFd5/a5diqI577MUfeHp
RRFIGhnK4O9IbcCVVkO3xoJKUsC4GzR29z4R+4NI44oE1d/Yr+HY75SJ0+NcdwLlN/5GuZzgCQtD
ClbkIW9QPkvt0GiBb+qeGXDLWlVU/XG6es2heIM2wVoEBZfSRX/00JV8OoDsnLjp2mRZUGbTiM0s
Pkz2MnPakIfTJliocQQx7ApGWGJjecZhnLRHypRQfmuTmFaQqVIFMrX/Cu0bcfOD864eggQiD2vu
1li3KDehJ3oBD4gO5/Qfx7EhgdRz++J1ZBYNwVA60VQj+xqmgetBQgS0Tokmho21kVat/kS2DZI1
B5dmLjLVZqLak+FppbgeZGj0Nnle1DWWrq24GTiuyIEQ39gqFiUM6RSH8SGk3eEIrd8cO4tnkt7O
Oghh8isUppjPAYvBfxSN6tKbNhafQqMcxilaXmikRDwaqHgtgyPqlsofUoNnAwgF93qNduWo/p3B
huGsGybHR+Q2yuPB+zz2fA5lH7J+QpUL6AGDKpTB1im+SxQD5MT0oiccVaaRnpbT57gwgFacvXIc
KZuMK7ffw7eEEPVRj+HyKGchV/3bVNahNd/zUc/RZJ7uKyqDok6rKGZoRPhwrr31Ksx+S/7r0fI1
ZWtW3jjgzjO7Bm3YTSa3QcvKJfuA6fmSf/x+aW6qPc6UauDnIWoyLI8YmmPtTJP3p2nmzpmVjwWD
x2MnSB1aLq8Jwwy9G3iZr23Pkay0ZOJ6JM2cHKTALnek3xNkJX8ABWMo/lIE/KchFb9D4ovrmDj5
ZzcdyEDU3z2Of17BzGkjeew1XOR8BvV3i4Sd1RlXM9w/QxsC3wrAGVOi6a4xHSx6fRTms1ZWadKE
ViGEQoOras6HHQb9Nv45NfUbgkia1sJb85eCHWImEhwUe3NLUKcOCZXS7Chp2CfQdfME4qaHQwj2
1+ns5o/GB9GWLzuHsdMq20SPkKf3FrMn0vM7Ka2iNq3xFau1A1f1hFORx3Q9+uRN+V6YFkSE9nFY
GuDw/96xkfuZXMVoWk5AcyGRngU6bapd1SRFolrseWfSYFw49QklzHDY5hLloxRBFr54hWkFtUR/
+48w+9H+S2SFI0DNfc3O+q1FF6IFjaHE6MmnY3CaQVa+x8aqeLPVjbezmzyxxt1VWn69ahJeFiuC
pqlVt8QviYJ8lvXiHpJioqrJDgLTbxh+ZE0h0f/rgpq5gkUVVIvMqwnFM1XmSNwiL4zwu7e0q8y3
XIRxOHr+sl1Q8T//ww/c9xcmTvPBFtSw2Qd9FAqKV4K94UiCr+W9aXnNM9Fk2K9DFzVOx3xKO2zm
mkFOwR5zLd1A53WXTPSOwl3782rO1XzqTtwx9PqJu0NsflPkbK4peGRyM16VuQJZBrdhxY3AdX63
QCT2DqV/7UvXoyX9GNQsDNXht/JmUGv9vYn0TNy8TwzgyytXse4+2s5q3ugSmDIo9GlqERdCinhs
cPfBUo2tfMcU9nNK53uosdb+mTB231JHrk/x9bXdoDVfIJcbnATZoVG7m/R8S4fF2Hben/jLkkB4
VhmnZh6rhHGBsFYQHuIweuPPcF421CMCt1np4NUAMCgDSjwwGkjLEIc5erDs5H7DG4bWur9Q4y02
SGmdx1/2kgz+sf//O46+SSrtedoy05cuBUktIdkn8JVVf1WdDtQ0QrA0JmVCaDnB2o3DeXYQC4qt
NwPURrIgogVosUbLyMKXmn40d5y5N59y+rPivx9y167xwSenv9kJi/qlVy5oqZyGwr7DB4E1xKCq
16GIQg0He2f58/67aq+7WBVzojVZdhhyCsqXsS1ahKVrSUNUSiJCos9LIVi9EYFCZsY8fKVdHGkZ
JmbgXSaTg+ModZlLImwy4AqW6D8TF7dvwym3NDMnsd+wamwXzrBnqHrtcIQXKjs+TPFicQwUnq0A
JPFHnT50oAQUidNhehPmMOR2IkUguP5wdJTBOqla6uXmGKLQEOdUP33Dzd1EikUisj2/LXy4v4Ow
WkxRqDN5PkyleFsRaVqgvp9CMYFCoijP92yX/BuBBvBl/NsFeuXg9+EFi6Y1mnXPMdgJivnVx2n/
Zjg0dyks5NowEWM5BQXOw+DpbT160zcnTyxwiFOMePWCbeAZL1MyEm7GxIuxxnR2SpbeRouwoB6P
yH9nbPaSqe4X/wect8NdgH5MZrfb1gQe9rdUe5ZjNIKuGAN694/SdX+BoSs8Kf4SpyLA9XqVPSGr
wO/In2dnWJQP7wwiBNLCZou8a8a99q+SCcYvGMfGuCiHc+xg2kw+yCLG3U2iH02vXCtzD9ejJr1y
3mk+DMlWKLU+PRYWe4kVo5fI/pd8CLiWawNzfWo115vcIAqIrwYUMaCCRQ2DpNTc/fmlmiXxg4IC
HPt8mNe+v6ZyUf5+A2kpctJ4Ifb0QOHn0GI8KC74RBH2u2Il90NkVHBsbChXI9ZO6SZ6b8bLW8RD
PYuZLuUNb59nVS/FxcYmE+kk0nVOuIMbwf0JrA/blAPo+mH8qUI08pjXafSbUhFezjxK5/nu4K5h
EeDpsbQFmNxhS8Jac31/Jny603js4bMHO29re1P2q9VVLXOC6/zwkx1ab90HA+H86bNixz/gCicA
LYxH3uAOCwHB7VVlvpRK9lx++266ot75OK+f2bAIDQQcn7dHkHrhzL/VhjyEh2wRTRpnJ6dCE5OT
9LfXABRTseuiOHh1AxbC7WWbsYTi0fGSrj0XP25OGP0LZ4cUPL5oDLHeeEJjxCohcmGt+HEgH8nL
DFnHBTWEzmcjhoWOH9dk1sR+53y7ioGuLZHIAsYggz49NMcoTUSp85z38OBM+S7hKAZVA876uEFR
w2QPu5gOK8RYboyXYF5pLOKfpAkfuGgRwv/uBHMhTiLKV8tvbb1opsVHBb+NRtjFzg3Xeou8vc59
LgMhyawfGMi8Q8Zptssvr3YkVTZYEvhGG142jZKSWU3wHM8Jm61aHLZ3hrKaugSs0kLqAFPPp/2e
l8sZJdCSjanopoU2HFbB0wrXWnHWI3KDOD5m1cQhQovBNyUtjabdrufS22/NpAc7I45Ki5QER1QB
onDgLFX9Nhq0xKiN+Q4JUsL06sEZ7PV4UUGGmBkJR954s+2vQSd7o2Cj6eIanRCkj1qXmdW2Whdb
1eNLYeoaXghU/NmQflmr3t8kEfDIR7AYamBpQaBzAfWkJGwnuF+qc8Ai7jdmL9un8FTOrdCFDLlS
+ImSGNboBhUZp7UCF/y16VfivClE+VFvpw5UtFVBESYPCtJCOyIxnIY8qjpoyEEJ/JGcZxXuRJ0m
OtV/YJdVX1EKSsPSf3OfhLtU2/qRxtQ7Kg/trhX9G/OYj2GtCNZUqkaYndwBwYV3QCpStxJcm0zG
uXROyGRrzCOS78BZu1rEeyPV7ZXf/hA5aESW34i4WFR+TZx2uKBzLFuBcISNLMGqMApz2et2jgKZ
G8vNaMvaKsVVQ5GG4ZZm4LTb/yb1CKlUB8ChjGf3CeR+I+9LzfMReMURpPtd2jJYGWK1WeNVo0JZ
CG+lTm4TWwlqUFah7G5RND1jE/Dj8Ybp/XlknFYOXazj0eDXyi0E1kkcgL8z++56eLahT+1WvE8a
JxPDSYzXpJQu6dwsTJXckjk4L7BoP+jja43YRb3a8gApbfXFm7j7crqJDjobCgRO/ihylNV/rhSg
esk4aWUoupi/DRjqU/hd5oqjfKKYpNDESBeKjEpLUCfBYw6z7PKw9G4I2qyIpdLPtEkYHnR43vAp
xRB1tR00wkWXr143TLtoPQUqqP9uMNLXqyvMb4/NTTdilWDtZ7CZIEXPt3RGU3QrbYIboMswHEu2
9AhDXf9aD3boeX8JOMpz2U3Tz7nYfv9qfzFZJQC605/1USU7xjb+CawZ39CTh+jn3SGE7zOJapLM
a+ClS45HCvyLn1fTbKT0zNC3778a3yn6tAzfK8HI1kUY9xTtb1J1ceXVWeKTHYKrJO8dwmtnXQWH
DgPXbCi2m3i1P176+pyuX2AjmAq/YYZDdf+eZ/aD3OHz+564iy0W2aWFM7/bxVageBs/97UieGcr
VpXEvFQnv1Xx62D9uxfGpsHVqo+GvbuFR8BNssr8HHa9RbqXptdUHTfkWv03MKzpeb6XMfpCvwu/
8R7ocbajZ5WAv6CupxE2zLpGeo6aGMB1EIeatBgHpafB6Ks7V3UEYgzacT12dVCw0cuJCRn/P+lW
7cHXDQMQJqjj8yecvqPzhZT+Ont0yeqpnMjqFlAwPLy8+HGGInmwJ6Ae43o3pg5I90ltsizFlDFQ
XtZNfltcudSbNtoGKPMlDa/tvQfcGbzHA588WVoSSjjribJRuQx2nFm9EOUNP9Ibrb0GgxjFFUCb
9h+zyI441EZKL0roujE2VfKdScxPc/SlCDlARGAyKv6QLHAIHlKH/UesYsWCUOBcKllLdPv8k83E
G4Fq5fUyE/el07PrWXe4m9WVqkqvfV1KAgo0NovTtnhYx3rZmVt7V8LEH7L5N5bsNrWDqgg+hk8K
TiuCTA6rsWc/hWjhB0pRG1DsWIpeivKTzThTHgUemrTrMNIqNAV23eNF0yEjC6MKeR7svjMmdHBm
mBouizFE/pYeUUg+titWX5QXMIWU+sDZrHb7TEHY7nwCVnvIkAv9WUqxn1d1f82QUMxGTHtqhS7y
URCv0RWqkcDJRVF2i3ulK4elvI0hjf24Sl/PkQV7EINPySPkMOLleQOfaOC4oV+j9IWTqCEQGucJ
3heYpO9kgjB2+7S687ZXVHKHUb1Xva7JspNwOp0fipX/M5Fkmc1EpDQNdIE2zxWpXBB52So7vdSz
/V3hazCEt7TAdjECJi0W0U62FVfcPCwCK5x1C45zKbTk++jaIpLGr+d6kM1pW5POC6zT87gwTgjt
xjpYU+186Ks66iCfvGVTE5aV6odXOOq71jwZx7zZXewfu4GyX8TcKUs9PgIayhL0nddtGo3gdM5f
TXM7QUP1aKFIbID2fTwNR1BZIAGFjuxtmuys9MUpb3/jKgdtoWapjm3JjQIpb9L3pDdMLLQs+5xL
fyyLIdYssXNG+azvyG2AieTrxBJWvYXAMqmzE6GVCOGj7sLcsagErQC7wT2eWnN5OMQ6yQFnQjnz
/VE89yMZQ5Sct2bRc/9nQqUmG++rzrsx5fURGVzRmTCuJBi8ApCH3uwJQO87MV/xQ3T0a4MTvLDJ
7Ocb63beYV+fEZVD98Osapbxwr72r4UclAN6oUm8sIPVYHh0lqyFdh+f4vcGs/jVzj5Udu2q90iO
u6NMJn4fnSRXj8M1GIjyiI3tPQCP0YecKLRB3Z4wiqImvKQtCA9EZEFtN8AB/eQmoANzKgRD55hV
PhyVpaPds5D8YOobQG1SY5jz6e3fWbAM3zF+2eWckWL9nnlAuoiAmUcZsIVhOAWjM285PafPum9w
XT8E1tDgc4MjbsamMa7D3apJl7gjVt7TCM+qYB/kh+jJ/V61104q0w/C8LsTPZsJ0GpudJkGzrO1
1ZDLdOmqhyn3Yf0g3H1MIs21mj30vcOkV30no8e/y71XmCdt+esuQHIpdPQlrnsGdj7qN3ykwOv/
UaQfWTF7qIbU/GndGNDS7xfcVS+ykI/TxMaO0U5lx+j6xUskYr7e3gK1GzUeTqGOXv7OdQ1ZS1dW
c+YO5GnVrvIEb++H/lcAeZlRT7GWy1aVMYEtGab9xw/5ggAxHbM2JcSNns7s9defExDqZXGN8gwp
BDB0yiwrh048HEndBDfIqkFpV7w+uih+ht0xdpGaTkPa0F0BwQSUNC0MHsYQ/eC1rPbFZTAW2+d4
0bLl5tjwFMTMCN9qvHctnRaV+sDGJzN5952c52Mj0sUAFtgsJmTwRhh429pUtJhUaWyugh9cTCDj
3p+ht3Ryh05xd5huqYt6pvvfwzdVLBjm7IuE5VOmVDHgq632sBGZrQw2lERWV88815VMFFKZ8KCx
8Ky42VbTsDgnSQEboWGtV6q63UV8BW2V3XPzKYsbGvn5fK00cItIvoBWKANggTBaYDot4gJpU6jJ
E9CbpVR4sGSs7M6zsZqoa7qpL8m47YEffg1/RJU419HEtG9GiSH91SHzkf4kvFRLC7i9phIeIEVM
P1ML/e/kbHJGrOIFe9giq5WwMo9JAhyGq1GLVPfPhY0F0vgLeMUvH/zpymak4Z0ra6Gacx4rXJMT
G/qYuSQcjr1fGtL8dcrLR5Ku7tgTg37+9GeAKdetWmibJ3LuvKWoidOdjGzvOlfT0CZGCv84QR5f
hVwv2aPRFp5/gZZZ5n4mmQOiqyIgb7Qzj159tThx7ju+8wE55prQMIAIkKmZyvNbL5u/iIVbBR9s
L+QW/Gl0y7nTGUfIust+EsmsEHSEBd/+scYxObqiiYEgT5AN+Mr0Vrl49/4pe3AGyQ9Bpx5+w0IJ
4BbApKIztbDAoX8H4oi45ivKpJSltHRNM3dlh7gcdremK04iMtuHjpp62Z37PsPUhnkOsMwH0EKg
MyW518BdvRLBo84sIwZd/M7oPB6U6B+m+7INm+Uuu6xPCf10gc5M2+JrntruV3NE2d90uh5GMzjX
eEQnxWVjvYxFBCM+uolu6xZaeG5+gMbznmW9lehKI1938oWLt8zG/u7SmuUG3Tz/BfL2t9BVzwmD
v+fegl90LOo1vVxzplAVpRcFQahqqbw/Mxuz0HUc3R6jQs+G2QvwVp5yVl3tcsQ79rEOIzptju4T
qXKd8iFFdTShR2VaTo0uifnj5SMdImdzBaDYC1x5Yturs9vGGUdzV+IIYUjeNVmraIsQhS1SpUD8
6rWeLo/qGd9kHdTYW8jd8D+hJRgqL8Awyfe/WDQJvEk0c4oDNPg8qGW/UAkQwqqME+BUjtkkGPZs
uMuoQlndIXsH63IDv7hiCyXsuGDK1Gqo7cnReGQ4W+CdIM+SaNOmdmqUSQB8VE5gdfSgyOyswrJX
MR619BAdDS1oiEchgO0aCihHg9t5JF9pFg5V5sCsWnxJEN2hMC1+p3I5lKsof3g7ih1annJOy9e4
CrMulYlaCpQIdzCbcWHCGxJ0K7rBMYmKAvB04g4Jm9MYbiL5bJJrUklxFg20mqklWhDPiTKx1fnw
PVwws1eonO4JwxdoHLhRaysFD6cqzgprUHaXzBPSS1b93d7qOvEmBtpUhut9qcEyHx66BRcCAl7N
ldtdo5m7LSQfRDk/dbO/xwEupiOHMCv5dijuF3sXHNy4j47Ha4AxeQi48B+J11Cp9NLtVV6uRaD8
q3sfiFfclW6WI5xXpiQAT88/Aw4UoDr7aYoa8sPSbpsOtzwzifPBUQn5zvj0w0Qse25oanYoZx+4
7Ey6NXw+N82MS5MrtBarGTfeNhAp5biU52qrrQbLizmyUvFJwn8tOSq/scHWpmty46hTNcY5EkAx
2O+vI+DTYxJJdS56wO+YGa9sDeuqeG53G3cLDXhkByQe/+XNgMO8kACgb6JCdgwe7J9VXmPkyNtr
SjYr5zc7aJi6oklNCizGKGCgVNW2kLtzBjJID2lgXaFKo7LuHj4KfR5feZWhE9CVFODzuA83T51s
mVH4F3CPlVhd98lc5arNIYU4Ci6IC0pq0+9anQDoHavRbROx0QswcPwlLUIC6yOKclxNcMHtf/Ex
EmqU4saGckPkzQLVrtbKZvLKPtwzKNrYvBPyaXsyBNLp9tnOZp4dEmaMOEiGoNGqwAbVFdlCCrhA
78OmtmyQXKf5mhAlbsoLvy3O7PE2MZTBdH67RWLp/F9Uvtvrloy178gVxYarwGRdX+JD79z5mokf
d8Sd+kQFMcsCYSNejhLtUVbLdiaFoPrDo8ZVN+HPxCEgeSMVWYECRaWHoaaC6ITwcFaHnTgvcS1I
nuuwpjt9UY/ATrLzssNimpfzzKKQCghVq4Vfe3zTY19wjq3UCqAXxEsk+H+GnROYF7hRBrKCNz80
7MTq34FxUuuozUERNoZwlVLxEZEtG6AOFw0FNmsY8vJMh/tG37i/a2Cc0H0067ZwyLv3K6HWrVIn
rNWY8Zj1j4akBvuajnuninHLacYQYK0ZdoSjZ877qZiEGNmqruUcO3HsWWHqvLFjY5Yd1F0Wrfpf
SfQFds72yE1AAtn6cBkUWI4Q0vO0p8c36opBDQ0HfJcGnHAXPWM1ZHsP6NUvlFwpy0Yr/4LSA1Nv
Sb/ESvqApes2F/4QpQ9D/QLoHgMwseY80OfS5pcD1RB5UyaM8WLjKoE/Oy+R6G0QXfhhE5NS091f
oSS9G9xZRvCVkn32Oo246bBCWhqG2camYdoxNQ8cdXcsLobDYH591ASHdVkZc+6aaULojvSDN2+4
PGNGKkBwImmQrZ4RPKsTnqWePfV8ZSUxdMwTKGRe6GgQ32hjZyk1AvzjaOMChHp+EI6L0W51IGCw
DT3g+72SvZsSQj0+A0prWrtabipWQRS02YZ8U/N9yUvhZW0eLdoFpCYI0wAY+nc5ZuySkBLAMslL
hMAjJSMqZzuAnXdeufZgOPvO2E/pZIuKAy/p0MDUWmC2FkxwP3veyfaHem6ART67wvMTKRmZpKA2
mAIcFn7NaxiRiK0zlg8pGvNfanwwPAqScIXTtIwB9DViYqWhhz65WKUeGXwk29hikhf/+/iPiBIO
e9HYFQCBk8zFnmN14qsjfMl24QlhJV56XIWrKyg3DRGlsiuyZxvqnbfS9qW8L4+CAbt+2xrpMgIJ
QIc3sJs/ida/dU1tcW2aHtnCrGI2jnTo6wqYZUTzCcrSG+gHOJxySOCIJIOSJ9bxerts5ztsvRUp
qfkxTJbhSUB4/k7tmF9HW7VlMwPAuxHrBF0ZmImyveVYsqNN7or4CAvPeKpIjnl/8M9zWSAcohYu
ZJaz6b5HxpgjO8B5GM78YJG+v9i7IDDDZNeqcFn6J1XpAlbvYQS5kqVqdrwuvtdwyt4ORESc19FL
E7sEdwC6feDYnDuBF9/P6iq8KG2YZP7pJ/VMSPNENZPatRjFQVD42wTj8nSFWVgRPDxY7AzFCEdI
ge1TXaOyEIejH9GskJriVPi4v5xUZRE7p1456WAoHhQmSwq88eyNcltV8yTf6cQfZxLQWMhnlenI
saWhvU83wTW0nkOyMHtrdQ0t5IZYqRA6utJF7CAe9WUbYPGgYlf3VKe/fOXpuHUOGBArclhz5Dfh
T+UwnuGkzlFExejM/emEOffZms2HYu35WoC6pS7F7zXrFLeovVamS6vP2esCGyXBzhY++1UlPRxF
cbAo9/CWK2mdH4uUtEPENLs+QsYV93RyOw0TDiWPz5RHfSP/tsXwoPctRDHrYX5ymP2HARIZ+oI3
gjHoqFiXDQdTjs570qMxZGE0Pjlvl1wRadWamKTXu/iSnJfx5PoVUtdM/6zGSTVZuFgJskj4uQc8
C9S1NmatCnVKKV8XlBUe1Z+engFksordXEmjopRCKAiWB1WPZyhPvycZX0xtff2WPpzL4ay+7/48
z6E+0H18eYJIBEWR7r7zsmp3eLtoM5GNgFrtP0fHlBpX6phA8qlPla7EH8Cx5HXuR/rvmDQvCBIq
gEKMod5jmpR6e4D9aSLJ+SoYIorROxTCxaa3ap/HsEcxVzvCcWaD88XCusm6KRaKY5tIF0mJb6a0
cjve2/JF8L1cncvbUewIAwYLVjGez7rYBwekVCnFbWWAaNkAqxlOG4hO0dwFD7OQeOrA/6TfaVPg
AgZVnjc7qh4ERR6xBs++Mb67BlmteekfAgvxKMpfMY3wyxuDHzu/v2c3HqEz9WxSO9ot5ixogVbk
eDWIIQyww+RCc9Fphy1ouUz/wES9v1o9ZOdv4WXJOE1Ax6n9CZs2RbUdz+4RKPWqntxL9K9vmVoC
CFUa8MztYxfvDJ0yZLiJQdkwdWsoWr/ldjAfC8tDYkWZkz5LO0xKRPXKNW2irNmcvLU0Xk11q5kG
UpZRxlMJO9OF4E2LOU8469ry3ldJo01UNRCwRhbttXgBX7Hyb1ZadegTcg6i58vPVVY0nSWZc4Js
Qk9BkV5Zof6YJBRGerW6NFTvgD3UR+HrHD1gsITJVpsWKCYI5kFHW7zhAHc39BBtZ2u+eKWIEH2j
Jc2ZKiVWZOp2DcMGVYHOzpHSMaudU2ltqLxo7O3Zq7Kh5HG7KRzCIYwMVyb291cXrYQ13BWfzYeL
cBrKJtrQ5pyVlUOaL66v7YrPq5CDt3kN+AndLFG0lBMfr/eBHNyKuNwwd+gRpFp6R/sWmX0UMPwB
jhCeEDc+40NVAXdBFNquVVQ1Zs4A/Oc9RNJYqJDHe6fm91nOaRnHThP+AMFm8TjpyYn1uW1CLV9T
Z/qrChXxyorozQm2Kj3camtQ2f22jM0uOuF3DBpW54HVtgdqp8ema509aLH0gCkAihav4JS5fPMQ
PXH4teQ65eeqA8eX11QYieeg6B3Uzimvwoqkp8SN8sTF4dvbcdpI+QcZ5qcEOWqZj1ZX5Y5YSRyH
IpilLO9DAqoN7CUsuclvXVx0YvIOAg/kyf3IwnHH8CPqcOEr40RfutVVK+vmXYcnqX0gNFqdXLHw
dogpZdeBxcC27MZgjfblkfJExGbEisVLpSETUPP9ceNGk5Vyh4Ny+bs3HQQflhQK1/C4rl4p9Md1
+y+iWyLZM26x/kqHpJYYElNGDiD/v1I8huvMtR05JM56N+wfgJmavKQ6DPe83gNXdSCiTTQSt7SK
fYIqPJg+dcWuOOAwDmjyiNo45nWVWWhv0dKLCtlM/19A8CwPEb5TY7lYtzFy0NrJMWUGwBhBLTfL
uDI41TFJVWOrtDek5Oqgo1/vzb8P/H051zN8MMqSykbQB+kkVpJD1IUqedXZ9jtM97gpBG7plSEg
+xLAEa1+FVO0NVr4E24BDJarRndTVIWcUPexlRHpbmNxAtAEtU/VMVhiiOWoxQ/2LehJ2U2Qzmwn
3kfn9PPQZPJ1WLO6CLFyx9kZSbelXuAm3TA7VUJNKUQeoS+Z2zGzU51CBv/tVVXaQT4+VwaOhb0F
07et5I/iwfBICrY9qgzmCbyvvOXbeVjoVivsY6eUb3FsGHirPW5wLqkeeoh36NNcxrw2c7OFl0ci
5vRG+xIgy+hqWTl0T1uE7GZkc5TqibokWjjMhPeGwjVO9rN54oUdlzP3xGjdlws7GzZ9DwP5r3Ki
R8IjToXKQVpNUHiOu7y///4CX0L4T9ozZnzMfbt99xKixI+5WkxS4lEpG2vH1rwYyYoDrsgqZwYD
8qRN1LeFKHLUgQDl4WwVvWAMGzYZJDj0Yi3CHjNKQc7gJCia1Q81UCthyG9jmEMpc/V50jotWa4g
rfPZPamB5p0ydsKty2Gu5jOoOdi96KFZvCIYhXb0l026cE3fhq1PUKqRpDz7osZFpZkbxb42GMm2
bvNHFf829WJH9OCoP92xYgVpaWIxYnfHF8ClrGgeqttk5yrfmm3sFEs4xHLSjHDQAIiz937sBL8I
gu5uJZDaFM//DnrjOX8gZu6WUotZsf8AcDm4UfQXucakMxpNXmiHDrUnSeg0BqpcvJiwpCFQ7DzT
3Y2UyAbkm3VZN8JH2YfBvcwLmHfK0ivDMAu1cHwAB2/4cpe9K8ShbCBb/i1MN0O/QGqDWpLYXzl4
APKyEFKssejMhBCMNR7h+FgHa9twwQjqQYD9KeP+LyMshReKyckidqJ5Gd0NKJL/RdUq8++D4xd3
jNl0wALlMIYvAU7fNkX6uf4kVtIOZcK0/Qol4oDMvugIRmGMMRzNcqrI2hjP0cEoMjmyMibVgXfE
4z7Wvxr0J6x8g5uuwEtyiOruGr1d+vUyZh7a1rk7eiIYlZl7wvDfAsjI9tRz41KdSLt/oJwB1k6M
SCJKEfNTLCeFQtKWJJKCRM1osAP2pzW59uqPlgLj2Nk6yMPEyF06y/Bhea+NvH412U0a1JlUafaT
VXS/xGlFHFANbr6BgHpvCNuFWH4F1ZPUtiViW5NFfJMnpBbpVSQGi5Df4xJEtxlbDIMVrccZd32d
L467U5yW8JObQW2olQZ60EOW/JJd96U9o+WZNlScXzxbGdAwUFVfd9FML3IxiMIOw1LHdlqL51xA
VHhkbt1/RaafYPZTmmBPM1dtyDjXJBu+ePmCMVoscE8RJI0kdaR0xFAmMizcrIuNWbkjE7odfCQT
fLsB3ZNe9Jeo2FvIK1ApKJ7jM9vihaPw0tfCep6RtAhEJ0Y25FclXsPpi9E9Eg2QIHZODvD7pmqe
TPo5mMJVaBOQUU3ZvOZ6ozqZGBzP5Yxy+lQ/yLUYQrVQ6UVPtfhiNZvEm5T0dsvctHYRXXducMfz
Hj24CwsSfrY4rDb3syoJKlNHdQXbxX0kUdWTpRjF9g3KPLRok+WhtjB8uUolEXBOuUNbiXN12yUY
JeRNpiaVPm9xsFuy19aeej1Gj8UKEJ0O1GDwvJaMLEnXdcDnpzA6d2b2iZCzG6tPKUXUgoqjsk+A
9gwziuJ3iktghEnLpT5nQf7KXDvl1wipEUydSvJSy/OKz/EfCUJePgvr77DVavDOnHR9LDOQHFUB
2tUHJQ763lJOSC+/o/D0eGAh/XxQbM03Jb0kLBEM1ZHoyd+mmmkeGJdKqttQ4x03eh0+6Z3IE8Ne
6Qgd4jMctvHlhGS4b0XrzhsE8kKqGVfHQmPq4/tfWC1MMltMmHeC69fFvQK59l5lXRuilv9GlUMx
E0HOZKnyRm69p33i5+CGEPfm9Xe0vTAh97eHtDp2ZVSG2iF8yi1JVeSOgPsdrlcuovct8C4L/L5l
flmYHv4NhJZsr0O6NWoM5WeJdo9HeLLjYkSlOu/wRxor1EhHe56b4IZohsFITs3ydeF7XZQPRDND
UIo8P+ZCXM/aRr5mA20teW+ml5DtJ2qJ5GEI+uhezDp8OboiMIeCBYaDkvLtPV1ZzqW8fKmVcwMY
293akQtQM/oeI5dDUL1ShhVouujLOgel5vUAzc9/l/Z3d2sbLZwpaohXEP8n0wsYgDiZUYuvc+aC
BbEz0Z/1f32WYwFeTH5K7kC74+U7ypMsT4rrcXeUrbNc0l51tIsBjpg6YlN+85m4gfjDZLd1Flaw
CWbn9kxb8RFgPovdAwLI+nsrwiJXwTYg2OfORX0iv1q4TiqLcecmvWH6+0bOQ6ipQnCFPKcRnGI3
yZI+Rt+oBAASWFROtrpk94k3WwBzJA6nMB2GRYBRGFNZRC/yV/P/Ir04DfH11E5/QMga8fRzJkwe
5s8OdiQni71btuEB0Cinw6JoPfC15uClqIT0QFvzgMHn0hP+2LLRGZzRqyiZ137AtL9VKvwAJDuu
f0p//cYbAkB2Hu8eFWvUQfaGTl4eYw2hCBkn7RDTpZPeP54F1YPlEzWhvpSKPtLuIqRBU6aBzeu9
uMTX48tGJvPuZ49lJWWVcrkOnizn1qFMaOahIziC/M/HeTU5/LC67I/FyfLN3CLsvKA0ADGLBBn+
kgxC9x1hREqglwKfK0Ra6b0ORHfr312PGvQ7o00tUpvAPv2Pe6IoaEtpXx3OADhCkpkgNU8xHFid
sImOLOhu+LRIRoCgLO1V96oXWtUBmhXIVFBEyPCU84PVaj00RtM2QSLiVOkJtWZAzpnFS2zFU7Yl
QXEAk23SOOiZxC4oe4BFYAZkSGWu8ocixSo9FmJnaV6XHWeh6S6env4yWpEC6K78wiTnBiA8eeX5
wj8iA0ZSKDABsJQLrk6cqCwITqAl3X1GzKIRu/83u0kbE7htnj0ZDR2lwcjVgI0tJdL0JDLYDMsW
z9F65fhMjCUofbKZUk1AMPZAtqGEO05XM/6Phx++9RNuAq88+iPvf+XFMSrgp9/EouayjtqSIfPE
tFS/vVDSMUNdlPs5JVFjgc6T5lOe2deln8ZRouTnogfNxIodQVju8aBcnJgtw134caiBNbibiozU
RLAKHolAWbJZTBd7K6L/YUtj53jMqltz5b7sTPTUhYQMebUB439GI2bYlhtj1oMrxXosYQFtjLwe
YZkHA1znjHz11pmIKARIAvo09YY2Kv2K9WniuLNsFv3nGgYuLQ+lsXs7LK6K2tan/gGT/GwEu422
59OO9n9IweTSOonW14RQ70ciyHylPmqwgHY+Ui99nlof3yny1c0dbifjQH3yJAVOZ8s4Kr/dA+av
yyRO6yg2D5AeyfjhsixnEL2EmqYNPdM8oUkknGrzY+av75ZA2mv0Jr/FxUJBfn8Fnk1DD22da5ZS
49oCCAPNLyO15uHC0jGZ3TCxsm7PSfgHD0dXmWIat8HVX2r0Y/oRK72tp94TwCscq8DnN9ZgNMNQ
ytFIdbu4ki1H2is154nFYEu31L42IzTk7P+YfZzABef+hZ1KoM7z7yZl5Iu/ddKgi2lH+SCuLMPw
+J1L+Hc0FJnR3mkQr3TYlOoPfWpOw4kyN0lw9d9CGIiv1fcCqt1uryXBSFjPmYRgR1ZVk9LugURh
vUA9myVwadECp+1rz3cCpUx+XlIra48CWC1nguIG79P9o7kNaM83xdROWsXlzVMajBrA9+gQtkXa
iBdvZQlgKA+wYgEBZa2IDH6bE0kJ8nNgC0HlV27/k00Uay32MkSYXmW2anvJi/YQWHVbdzXy2ojg
vwfHfAnDW9KUFA+OG0vV7dWwlZb2Vy4ElEFLUmn+aK71NRWpXq5DyBBiEWmfbbSFyTU8OjrKFTFm
84E4Af3M1ak9VRNnWleWUOsNmqa74L7kZvRkdkg6VuU0mdreOApekNSs9wMC4gE8+bdgCzWZch3Q
gcZocYm+oFItjbzbRE7LiUoqconFkgQTzpSTLnQYZbVYVbChBB/jMxUeTvZrP38YPfC5Wl3lLC4l
H9psng/WCjYeNxkLg8R/rHDVIdugkDXkI2PhlO59bjE0LkpBPVCD3JzRBP552RoNT2kr1rQjUAZN
CzEwX2ZIGRtUqIoVcT3sPzpmJIgYkKFRSMFPE/C0VOZdzK52jc6FAlx7kSbnudfk8bq6Qzalh6lS
APaYWaeHJo6WawGzbEG7OsK8u1Nq1s29ecVkMmmDRfCl+c3z5iV8u56RU5O5lERLYXGmL4biSzzp
anSd65GitlXO5yLgJWZtKqlHufN2T7UqIRU3zuGxepZmGnhLnC3C77k19ZET+mfiRUdk6h3LbPaD
Ub9gPYFV/0At3hqRO1sW4HMxVFOCJsPfwzhX2mV9fwh3khF1jglcE5BmqIE2zZkV0Rg/ULs/m5Kk
AIEZvJTdSl7MlJsWmFv9Y3t3ZD3NQ+P8vl2xDkX63qTmg01AchoQW7vVaQy2q7F3KzHntE+hui7e
Llm5kURZTKVE3udTAXyPu7QU24Q3u1GueEz5dmFNBvTbgV78tB1R09+8IuQiya5uC7KUwo8cYfaF
KGI+PzncUvZNj28N5Jbi5E4vgJy+lkGPMmVX75xQGzIoSxm8KQmTbZWg/RomjC+RLVzNY2Hg5wyq
ORtwk/JDMvdALM0cYN0datCd7HXhWq0iAtpEYAEPCc+cBsjVVADRR35LSEXzUrdWDHMUfQLgsfPg
ca/2oxP+5h+MGVvobV2l85suTDaWPraf+Hp9qQZXVj4FJJ1twNmIMs9iTJJFbGiVyA1/YrxDbR73
acX7U8y7bCEfv3BYMrCWyO/NacW/yqhNxihe/8+/VruyA2mink+gNk/uyW5I6RNWq5o1rybnUhtd
Op92p6rqJ9q0yVGrMCvQkwx/w28rmLXB1PMoCpQA3RlBxzCpRG/BACLXC/6HAA/TmWGmavEcmvAw
m6+JJiOXFWHcquaF7MUQFQ6yBvbKVf+Oofvrr2yLmQyiFWaqemSwgqTSIq90idWWw0WDNJLiZXFw
xnNswDpV7r9XPioYWDqq0JhYE3uOSe1oITRSvjjnoEM+BTnCL7BM/MYHkN/WEolTIjZvEp142zd8
Zq0pIir5MgpClhEa6fksJf9vex3CArzCsKmjfW6sToSiGlufSPHaRGKKGpip5EoM0ILcDw6uaS8P
FM2SxX4JKZUMDCFh2tDoWohofoXQPFweGo8ikn1oAkWj0nCqo6ShcQnj7gXopQKHtIRxAHu+Dx/x
jnbTFNv03XIn5KssgJJzcasuRRyL9ggHwU0Owkgzimq02xBQOdnkQho4cLLEh6Vy5bZvsu/j4U4c
I36Rh/dpC2ZYmhhe5NpECKWIr7EQPlto4oMfMDnTplu6HKG93c9rJpJEoUBqOvBQEdwuQqWhSGF7
uXMXIy3RBaECVPrUpE7nR7QifP0oZBnZEy6WnDMPrrTy0yFFXao2a7AvB1PqmevAadVSzmmxev3/
d8v5Io3PWhx0k9K/QpvsQLxL1Wq/zZ5pCYFPDncBhgRE8R45S4u3icRGpszdF83zVlmW5N4s9yO9
XgJdGdxx9ywPM31BozMD2Ckjt3h4zEvf2JyWX+/c50EKEsbJaY2qilcsM0fst89pWse8iVvvQv15
NOq+suv0E8mpT1PpK7YI4d3BDsZ7ps0sTCHPMs2mlsZOnzysyoDHULiXtNE+Pf7zb2G8ilARGIf+
6rQV9kYEfu5XlrTy1J98WqnCxPwEhdLkLEAbSBQQvN5AfEUdAAw3A9ZH4n9boPZJwVqc7nHCZK+X
giumiLkJnKAn+h+NEgFOin/1H+Vr2sVI+pynKMVKYtd2fwQwYZN+xhZw1FR0MEnHgp5c26cnQfQ/
+GNllXXTn0CUtxo5hj9Sgy9iGDCj/oh26Q99oOeRcoJEYyFF82roAMVwZHO+rjbHXU0bCh9wujsi
Zg8Hord8U1SeXe9kdGAe0eWmDHIPSe11nwmnVqi1cQVfGSgyMZeZebHMelJ7dvAB6SGN9S7XxWkA
X65lduT6ceOW4EF0mZVt53JmWI7CGgvAeshiytFtUXYAz2qkF1W4sNZ68ysCJ8RRN1DFaHdo3hEJ
PL36jiIr2IRxSkT2KIXRDdQFi6u6tVINilgO9SwTh7EQyjE6zEvbj2a+RK83I6MnmQx1O320AkAE
iSDQ9MQYl4f3ciCz115H8ozWnvJHp8I1z1VwSIguXxbOD2v1secUmQ39Hj86WODJcJw3YMZi7fc5
tAUUT/oRxDAq1/XEtrW2vwqxYDik+nn3azZNY5p3NeGZ6ggf3CCT5tlrr+BevWXE1jU724dFUYbg
DQfAVw/Meg+UwOgsQwA+7nnvzU/WR3vfgbWmVKRiR10rpNrfUmhCpkn0oa7khV/6lf2ucUmU5i4r
lmVA6Vd9YI71oc8LsDdEEVruQ2IBA/8mlDRCa2io521rzHzrIE+H5bgbTW2pP5048bQPb/L88amD
iyY0GwQDxGx+IG9dB1HxXbkKKomS8c44+8ZKj0cmqOh1ROrgbBj2G7t09/PIvXiU/5RLZuAvCs1D
ThEDEEQz8V8WatbXAqIZPXwxNWX04HqzJCkSumNpKJ6B5K6aMCiNgDNMayqPCgN3PK25UKqVo5TC
0FwM9Ngnp6CgWUvRL419E0ra6ydAirI3SdDXSxNXXM0dKnIC8LWDep8EKVbQcrLuG5xu6n5pJbgT
/VjUii+cTKrMkgmD8m7SP4Nq8bEdXu9I3Lv4iuMlJAV4zi4LnCtW2pVfYA7YGxa0QpnRHxzhe++M
MRmW70H6Jue8kwct/q5bq5SRhcCUibinmcptEryrjMA9VslMqYxIA+yCSqZ/4prSvHVbv/mDuyCQ
/uOyNzTc63CL8IXjDKgwHbXq2ptDVF/8Z4GHR5emPEjruZRQ2ndckr3tQUbe1en6pL+Kw6Rxxn0Z
wqZbgeI65BHFTDqhqfMmDu5Hxm4r0Zrkxznj1vk88cQddjpv/YEH69omcWgR/58jBiMmdyYVfKUy
qF7Tjc913f60k4DQL99sriG+9HKrIWBg68HEI80A9oft4jwibSwz8PnqVbMnXW6fGgny1mjiqAsZ
7GA6VvYvqCYybYqpJGDgY7wYMSZljF0xVtS8YgQqVIkSqJij082OVoYrduLlTI8ytYN/KhQB8b8j
GHAf1a5fBw0Iq0KBsoExToS5esQne4afxykdjEz0bEtSrdKacU8m4lMYQEWmWDE1Bp3172n/OwaA
8OLFTl9hXjuLvFFYaCU/1BLp9jO/1Rg1COmHlWTeIPcN1y8YPceqtwm5urpbgKlF4K4iiXGAPRLB
gvYVWcRhN2kg/nEIKhv7ableI00I9eLkcnzQQWr0unwGIS1SG7hp3KkSHdQ9Jy1ciP8lD/RlCVt3
F9IU7G24guLilLDXQirBxC19txDj5cXiC5fc12R8fQh2mtOHWzb/pud8AyCQtgVmzmwCcp9KPN1e
A3rwdPfiD5EV++Cv2b3/846AObpb/RNGWg9vz6UHddoghBBJb79ubvMi4mVJbNFhcaI2Nz1TXQEH
UHRkImK2P0eF/7f8zt8vjSDwthYk4f9IGS3ycdFr++o2dzO+Yc5VVQOm15+Zg2/18bfR8PmuOrFq
fU6CsjpgrALI+iktole5XAPA8zDeX8MrNiajlIjArJ530VRWcLSXQ+uQyoe+9xJe744FIvpEp1mO
N7MFhEWDoGw4j0l7jrOfhhkQ1ejthi+xW7KwSybzer47QsHa/nLM+THqILAQqwTC/Qwaag8cRnWb
3kIRM46fA9bZ9XMP6wEgJCgGddDolIUkslsj8XJFf5pDWQ4KQQnpu5tJKt0gVULGnmWIOnp6ysou
Kc/rpxKkKOcZu4ygLVPDk0PJl6ySpIpc3a6NELXEXH3vPpE2K0GP6QESYXVcEBdve+u8JwvIfDlx
oSat5jyOcAtBTD3+EOyS9YtT9TnMAe/2Cz+qvlEABjQ9clOsd5pOAITu4pxFcgk9YLtuKlquS9j+
my3mbNR/N8els2mTkVIkhDI6E7pBWBug7e9EsKYoBBDEltvU5ypfMDolXi0lSeTg6Hx3yLnL7q9t
wckedDqSqRfqv0ktvt8TaglVEJDyIriG+X2E3ctOIBF7+xMfcXzE8IE2gpqTfU9gZhNuigyq4ecA
2SeRfJScy6wLeIoFbwPdSqiU7+HAkbmC1l9XnBMDNrRuZNL3yHTrR/RZ0bimTP+chQKuD+7c/nPv
fz0Xj1ZM3I4Iy6qYitHpX8le+R7sL46sXlnyjvy2ETSbvLRyzi/1JHtTuzB62MNeQLwICnoOVJ/S
01RGUNkBjDgoD5Yh+AttP4fy87NdUU2m8s/09E/ytFOXixXx+2yvxOjn2JwYUjmmXiw3OBkSiOgA
oyVhQU9VtMy9B3EfxJA2YKyvNqATHxQFAj8ZMfhjAquBw+6IeYR8ShQs5e2ej272X3pLvvgyjF0x
JZgOTSM6ygw5MMGfl/2M83ODFYwryNgecJAPqizMptODe8/mHvl3iPBVXmharGP2Pe4OsvZOX3kP
qN/YdeEAfox84agxp6eu5JUoDSj8YrAkgKPa+NRGyGSb0uxS3s/3qBlGOwguYS5H6RXK1ByN0sv2
p9SouQKIrR5T5F8BGieXplxspA96HVpO/e7omGiHcbgq2sTrFRzT5bDRval8ZPgk4OlrBJPImigL
e4TI90W4/JdAZn92WdqAj7t4bEvI1xTOboKbb6V9eLT3YSDJxbz57azsPR/qqo4OnpBprCLSKuQ/
5sJISdjg3CMm3WRsFclwWTS2zdZI4+ooW3wyruCKbDtVQPUlyqXYkyixyAwzCDXxjAdFSf+8XBLH
gczKqc8LgnTnxoNU5Y9U8pJmo2aA9IyCE47vapvlbOEn95fdXv6JeOsdU7dMQYhTWlfti7+ciNiv
CyN+PtzZmr2zYzD8KtxkcTTb/d1vkfDAAdxz9rzbrLvbmm/VpITlWj8lReA2pCa14TVA0xhbSlq9
4DilM8S9/v9AjnBm8xINIJhyFOTOZ1CY0Mo8lywmwpddnuqpAN32Zb6e09u5eCGnUEKvB9urcGNB
s/HDVGPMsLBDGBDdmMT7s9BjreqG3Emke4DzWErV2CAi9+oAujolvaYA2BkqyoxzwD+wog2JTLd0
BimIwHgc0XhrUksrtTq8n6b2FWml4jdax4XZMKDBdHrPY2F/08oRmHSzrYCSNouwYSaS1bIhawVv
QV3cYUCYGb5YX+lbo+3WUhHNdkReW0RMMD04sqj3XVijcnkerUY09mNni3x5W6gKhXXqsHNGOG+f
rXaYnSCUi/VVdalh+S+reL7WljRY8AAk1NyKlrzRkk/EDiupyJsR9z4G0U41GfgE279sSLRtPPtg
B8JSt1hNS2E3RwGKmRoib7SoQ4Hvs3MWSTVO6K6vEo819F9vpoeBp7JY5V5yv7DEzkuxkW0knXiF
4LH69AQXslNXjc0QKsPLwEqVLEUyv17X2g2PsCRi7g3CFc/NgFvd2XmV8POoH2lW2IsesImhO08P
nADgpZko2i6na5y26lcpGeD6lq3/s2znCYxYHLbN/M1sEogmDPm6QKoWhLoBK/HbnxLkbYEFH7hs
2d898EH6TaH4Tj4v8Khow2iyogVj3Je3gcBaau0rJgOoA3WDU8rCdMdU3OL+42vzQry/qJu4p7Wr
uSoZj+uQYDynEj7gwmjfmSlQOYPi3Tweaom6OHqtHVyw3mS84CxKRwY39kEACAk7BGe4VbWPnFt8
AuDo4x2udsZwQfDfD9isVKq2gFYSnYma+UZKChtCYCpeDO8/3ImiBcf+ph9qewIK/pT2k2tKYAub
4Febr9iS74Mhkf6vbOsahE9eCd+zYGFITPYhkvXaFYvny+CBwEaBSsSjlIiOnJZBRcrpcF7BwBQm
BwSVNNjGQSVzrpw7Bz1SlOGJoMcyjdEMEoKOSHNwc6cwYLOVzkc6A77+zlqqypPyHhyPKQBspika
euYVljx42tQ4UV8wDjk4oYvd10AT76HcbnNXghYliX7fOyT6jhEIkTMSU16s2++WdE8jfvRDOQB8
rTE+12GfwSsnuM1ThwC9jRu14pWciVGJitVOgpxin1uKHLc/VXgrWCPavK1qze1M2MY2BebdZey8
g7KRymv9B0t/YPPMh6IQRYc/b2ySxTjuZItS5kWmTznZMpDh2CUCfw6/iJ6RscjiLDKxLXd2gv/C
1VrUUwwts+KJ4HA70bg3mdRWOcJ00GRPQTM5bpem35/Dc5aG3tTXVPI4+OQlUCjX/su+/KwWFLgC
Wsb2YIuL1ZkCF+0sNVE6XDb4RCZ2np6LOkylqTExA0aO3VDyEkkFEUvLnsYEN4uVKo5xFkbC9X8j
RIPENGP0ihPchWLIH3PMAuLAbg9898pLp2nEgaS1iJ65BZ3VaedVvNnfU+j/zQ4uhKDgJl3I9iHg
oWoHY+WAkMo7B8XN2FynZgdxOrX0k2/6nSfqD/dnyuzw3qMb6q8Nd3GuVQYHTyV+YBmJiByLzqIS
/icydwV4Il0B5zmGgKcuUv4o0+EM4u0GfrIQC1w3l/9p44VjmArv8JVXvwLevrrBPPrxnvX4axRx
g+70Z1+ljooxpKHeY/PC9F92RTF7wi/idKMh/uOPmNVvaBrtl6Ywn/MDBOIwefBmKEbeZBZ7TjKF
rs7T7fmCyCJVU+0j6wGdYJEiJUScQszDgrhtGVpXFKQ0EcE7CYR0Y4ohD4UP507WLaL/EFaMMxUq
G8ILunbCRQDEpF+XSTGOMDpmFoef3nov0Yl2YwWBkAx19obPE4EW1Yo3ZmaeKjjDuntIynfWcv7J
6rf+WBqPjim6SvUCN6MzA4st4L0B+n2TRRaZIpdSCGy6ADtdSG4KjeqO7JlCKKKkHv8sapleSFG1
Efnk3bZSAog9xw/VK90MNnVJYDiAU12ogHsUn5Lk1OB02yQ9kNrpPHVfuIeuy93Y/uIFe4WSe/5c
37DdbD/CXGb1sm6AnWFTegXbnAcTR5hAuzyfkPmNBY83blENGvCXRIGbr3RUFb30e8SnotwOUBHF
6+Y/ZWajyZkQCkFY9DKJKufREpDR7plOcAqifR8usH1g4UtOJAUJgwXlZy53pLUrRKFRn0XMLZxI
uMvAK8NSJeok9NM+NrwGH17O7yFAoBmJrJ7/35KsFa2hTaMjDGUVxhHZJ+MzZ8Z/W682jJRDuEa9
o0IrvKOl1njR3LEGQXl6lllFRcSCsnIw2gUlAHiV8hTwh5jedhC9kVBALgUn8qoaCwboYGbV6jjs
Ftw9vBFgzx4oHF3qAGx3HbphFuu3cyIT2TOJef8/6ePO3hWUOVPP0tnCTrbfHeSWZOJh1z9evVDz
qFgwrre39chOThl6w2qeDJUDzxeZY9JgvYWhGLUmvJrlVyW4fyrNAUAbF6wu89CkRWuTYGcaAYeh
a+8zDwsPHD2Mcl92rbk0m5PMZB0YcQM5V2EmF1864/Rj+q+2Ac0K05bsD6H3XeIr3OJ715+TemAY
BDTRRnDStFD4p5iG3faGebcX7E3/tavM7YOXh+hEs8d6Eix4bKwCDFaElCs8YMlRRPfnORKBMwY2
nltPOcvkFANz+NsuuBICQreemUW82ZEH0I2t1O6tiT/wBWQKIsyTML81SIDt/I2U5mAYKM/1qIlF
XXmW7G93wojmoDWA5Y/eaHXfXZj6kKA8USV6z9he2GOqsNYjo4sJTYF3LoTpWlakyUXBm/BfUNey
AApNTUaAEBLc23MOCsXauy2LZ7gRGMXmBiAqYKXeTGYKoGERNNPp8vg59gDPtQcjUrb1elPq9R6g
6F2emoxQWjxow3KfX2JfDLc86Ao09Yj3vnf3cIUGdpSnAA2UUK0fYHGmOVVJKXMRNkigEuOu96aK
4bSQhZZQVzuDqIekxGTFMaJJsC/MHLXbBh6viDp4bklt/GziQ5HHn5cqIe+dfYzuEUSSbK02YaKy
6kns5lSDohdcDwdRaj9+2kQz/b/O5E4AVxhFR9D7sEny0abVTrxgfCmiECG7eqslULK6b48aVb9/
G2Lmx38lWRSuMbknD4cqZeNk2JtnwNKeo2ePPpHG6KrZLMkZZFytj57JO4ItgGNThcDwDv5sRAa0
PBoWoYNrsnKPfLsCYbk4BCJnRii9QtCvHVbKs9A0g222RjmS1vnGDpXwY4Q7i/0suQHXuND9Oufl
YwQlvc2giu7gjhzs/LAhrGFc5u+4KAG0cHBdmX3Q82tsSgVzAmSNUav/GvOryjTyG21pWKGOIOKR
Bv9L02sqgE+3FEcXvP9ttJwMST5b9ksBxuc0VUk2vR7zvpY9ijIP+JJyBVFstIsBMM80kyFm7UdW
DAm0eeAdVY+X9kVvaY6FrU1fVpQBI88gEQ/1+Ltsgo4AwHyJDCxefUzoy/tuvHgUZNPDuQSLuB4g
XC/ALAWDypVfhmxcRWbxNK63rnlrN4uIPyVogndL3ac/CtcdoNeiy7T9oM65aWxVjuoo/15bmHfC
3DMWM2J082EdG6oULJXgKBoAu51ZsF9zRnpQuL/6IW6lWQkEB7OIGxy2VzRAu7IJXh9X186M5SMK
g5gFUNgkNA3VH9I1Xuy+ZSAwtsY+WJ6xMRs5V8EN+LsOEcCAsZ1pGliX76TMH5qfV4hmxivPJ5eX
17kfmgUzV7V36MYL1qHNt9iRfNFwjAwTFysbcEkG0dKSs5IPChlNzXCBlGI4OJe7EAiKAQCZtFt7
z4rWB6sNJChJdI7tsc+O6slJEubOJUiE3/xZnPL7uYtiroZZv1bWpwvTEb46/23fQPIOx62P80YE
S9Be7UkFM62eOe4QBkrDDbW+W7bZqYFpBfWEacmc9IBg9g+KxGUabB0OCjkPGNKJycIDyQmSQGmp
PodgLFyuUPv0fzic5j5SI1LvYq31yhbTohUwfgkePU0hWuQDHhSotB7+FGf831ff0H6Dya814cN7
BeDJu47P7OpH95BhuJnvA9EBztKLrUJne0jtKvUyLhhI2OVWP19yBb6qgGLazskHP/AJd+P7B42v
kZx4KTp72ux0c0k9Oxv+hvJyFT3BGD7ItshnJ+3J0yZ++rcWvU6dX77I7biArdzgde1p8QgJDrc5
AWF/0GthfcXlHHDru0pFVju4jKfZCxTK9t6qAGUJXe4UpyrG2U37KtSqidv94zWuHfOwRnTtMkHF
YC2cebmxiwUPeu4OphuBqreuEgQsYkrIUpewOSJgZf305CanEJOI/4UAdOnnQXTjigJUMx9uozlT
VStsCdyF8LT4dYSXzeuPfpm8VVVKxTzM3TcTwvHNCxh4Da5eYL3TZV0kG/aGR1aezJVeeRJBJ8be
YIqYkYK31MaRRtQ8A/en4y5ex9uRWCWAZOSBgpnHLuszX64BApHNI7RRQv7NFoBcL5d6br/5W67L
qsgZuFMVLT4NyzjbKDEOUv4LmXauBYehGbiB1SSzcdGbDEtWPndRJWQRglAnE/YomZExt+6WD8G5
SMUMk6HPlX1jDtNEeZeu6F/dD/Y59ybffSW0hRhvl5s6/8UMGQqiaYcHd7BUCFri2cQBLJF33n+0
fuJKF8GYRtzWHRZxK7RkUVGxib40pzvhKEur5ETSKmS2ZXGiOadUyygJ1ottyEHKOJQYX9KAdiVs
gvNavpxvI8cFM0ruFYhYOS3Up4DYY5xFBUGLtw/UzgFRgtRVWpALjLho+Ls9tZbJiOR5TZZns+sz
h5xtRQT/UhzC7h04kdzLMxeEwZQidZEruOS09HweJvD3heW/czsKGXjfWXTt7cyHcx9DhnivqFIz
vHpyLsKriuq8IILxYG2MkjhhMTKXXW/Z8aO2u47mthH/QAsy6hb5UZT1CXo1dNwARvzIovrxoR5I
CBT3i4FrRoFg1xQGdo7yhq4z9EKMATP/abuo3zsK9z7iTJsr2uOH4c57RosXGrlMpS8FcC7RPDMB
oS0Ef1DPTIpKoPYPbE3LZA8J0Y6spJkGHWfeWvwDBoevCYU4sBsxEiduFCnSYIngpeHbc29yzdZn
cmT2+o4szpZL0DWXUrWZkmJ8jnNfqJwHrjeHECWgjsPQiTbZohq7yKqFN4BYYwyPs7KqVjhWsW9k
elaHVOclcVTvcjPMTEvYSfuSy5pzI0omY8PzOgLizBlfvwWHbrbsQGV+EOl4w3JzEhlYkLQAbeeb
9BIQ5lyuO9R8ukEaHk1nvYTt6Dt2Wv5aL2h9RY+SQfnNldCahOmL5qlqd3+GDBJNsisBvq6TFmCB
GIR7fSuNdNai0bJlPYINtBAuoal2d4wSaK+FCFVpGJhUheJ+pyrVKSIi25MoceoPSM3QSem26zBH
btvjuoo/6RVzJB71TYf8WtJkRx90X1oQscUPA+jxNgoulBQmNIyJIBWke9fB84vuKsopoYbDiY8b
xT/P+iXi/dPcmZ/B0QqJ/013B0yPb8ZIP+zjB/oYzbg2grYwDVT8Xp5Rihy6bnIjxX2QdWFrZX2p
kHfHE++5Q5KqEqhEwYMH/RV82lwJLXDYoNJnFDqi6WLSqZ6JjYQ5cXCXdmokQSJ/6i0B1qtqu3wA
H96fGhMwtAXBYc4jqdze1iFClBK3olR9gIn8IQyf0h181+eaH7VDxROCTe5jPFN92Aur7lWxUbv5
yeWerV2d5M12JFlkFTHhI/wrCYtgN7HzB6bEFVQEdyrGpmkWmPJrHTjSvmRHMaHV6qSgScvkHDQM
x63p5GxflhWzFMwThCQzmZNgjdGvfDz9NdgSAceoiQ7G3JIFm91YEoGx062E27fhAA/1DTDYH3cI
8dGI2zj2U10UFC+FCO6KTXqEcqO9zVqbvPQUxJXraKOyxgGNhjw/vyZBey9l4NQ92FreQZP0RBeW
arut78DVBZqO1Y4NYv9Cx/4IARV6PxObZHo4bblB4IzKF1PgR/57Q/LUIS6gtOcZS8KTZSHenWfK
HEWwi1TTBTHhIeHjDa3rmtCUQVzjZZCn0CyI+ZzWGIINR/Z1/b/PHg/KbpWu9gibjcXpDWhd9Qhc
5X5maDZ05a0MkJaS4F2GrHkEyUQX6Ff7l8NOJCkgZX6rfxJ2m9P5IMH7KmpXootODG6LYUi+XPQD
WQXkme7t2juELnjbxMWqhnnllh/z2y28+iygOyrXBHiLzNq7swsC2wWRs1UIFevrQCmbjZFC3IgS
2AqXC5G/olm0j/4uYp/6MozIG5hLgDKVBl0C/ez21lrnrSKp98w/257BtRiLu83WzueJapg1VYHD
dT1psHC4XfjMnCPlRSsK7QYBcW8ynnzx0J3c0XZ+03NIYxD245kzGGA+CgGViRotffWziYT4C2Bq
xn12gyRWg1/syGiKCRJf4U7fstGlJDSD6VvSz2nPyTHUFfDfAumX68G3aJdQzLVzZQxfcl4CR0on
CspE50D2KxqGReDhTbSOMr903c98njO+haz29yzR0HzuYRtte2vKfUeT1NQCghNnVkU+69Y2ZX2K
FZl6B9f6y1ftTKQTZsSc5RIz+ckjKg89boaCXNnTR/K5H+IdATIjDc6bPWRe/hSeSQwMLalaK90B
NCG2s3gxm8J1HHkqcLjY2nsUUgmwaHNFwlkIEnYhLNvxMVT2ERU6bW+Xz2sayfR47GSV5Vwv92xt
2UPNqd6dbkxyK076hB56rD8Ka/q1CtgXPNnyc0BgtMwezrtR8d/lWtTVQSgLwj8siP+do6bNDxJn
gBuuiVFCKMniCiEt3WV4vzW+t4W7OaxEe0g2lHbxT4/HVrpy6iSAP4bLqYqmDA+xqptpE1nhBD9t
fH2PncC2tqK/jRLVM7Nu9HfrJ+VK6Gig5/+k7h4QyBjsh8eR8JvSiF7464NTxCsM/idn65dFOEyu
d6Rq70W1MmqjSCnZeg9maSh1kPeULsZHXG0y1ppU/nCtZy2ixET6hFHdW61xt6eS8fB0a1oy4tMT
FW52S0mq+FnO5+B3wE/9cuUXQ+sAh6mWEAGRmRDMCXAjl/4QzBL/yQ93jdtZHH5Qz+HTHBSS97zK
h9BdYIDHyzWrnKVofYbesUe3yuZ3BhlJAX88hT+w8PS67+VzNEc/eAjaXnVfNM6mBRCHf7sS4NmJ
onXdaM8JhfDlS1lrop1KK9ckJJ9XUdrUHZKvMNXuFI6MMA0Yla3WaGUZtiGK2YYd/4Q0vlQ8TKJW
eqoGqoLs4uj7PudB+nwAaLHSjh0lOGQP0r1nXZAznhESM03afOGYMR7chUcvyBM0gN5nlzoVKX1q
LI6Lnk9CCgmtFn5/FQtkDT80c9AZCIst2DuTx9gGXvMPd4CB3yAl/rqBhN1sQ6YJFUeJV7dXpYTX
9eVL4kDJpOhK1RHGHNWna9v1au5l6Yy3tF4WZSHtDufsgH+0cwbQTXhK5g+50m4WQ/G7v+Z0dmDZ
hBb4S1sm46bTLURaK5V8DiJX/o2ybd4B+9lklylwmVpQZy5SDNslks/pMahZRAXcGqb+/bQi7BRN
EtS84/8O5LJzCtXzMzbJzCV+B0XNWBBzWfhv6YmsVhwdjrBNtZSrhtALY8BLrnPkK98NIl3mb16w
lxJjiJtJKnq84Px7NqRnFJBwr708fw66OFu1m+7I6nGuneZz7oHhUVORIzLlpIOLSuyu+l4a8YL5
H45CpNJ6iMism0Ww9Cq+v9Ob+1bONFubTHUxnM9KOTPc72xIytx/APs3HEPSr4XJGDOkaH11UOYG
JpJkI113XgzDDNwJ5o3ITDu/gWZmBqlvJhIhMSZVVhBjvs64ZyPPSNSdIzbhVQ2eGh0CwU5ACgS4
rjI3QmGhOprozH8ejvKJnYvMJ5uhkbyoAziO8uCCl6tTYS3NJ7jWzpA97Yk8Zhpkc7lFh9S6JaZ5
SNLA84G6/KUGpO+WGScVWvDo7+wcNvyeYkWQA5ihooBJblr7fpRw6Om5ZDzsa85dvjIww8F40hLH
0Zt4nye/ou43cv7r7GyE3MULBaNqIud7bpNrA82FdDkuyB3KhDyS7eiLGb0rmTDQ6ClThuCiO8XM
mVxcgvnwFm/Iga1D2Bt9XooauoTM3bFqs6yji1Jw16/TzfXPi24uAL1WnFBj8C/rr/p+29fu9xhe
I42nmsWlROZSCVTXhd1zStWGKhJlqWn/0nCXZvw+4IZb1JumbJvefaWz4dXgAayxeuhDayn3Gl9X
6syj/aGnN1BtIFiehVsgNfDJR3o1ZD4sxffe3bftlI94OBe1/nemPlmAqalTtFGD9Ra8DXiWdVUQ
g5JeRlJZVLy38AbnpmEkRvY/rmc0wLYi9qBUb6KFPFsugWPV1IPcN/y/Tk4H3blbSvdget0SpSQV
B0yutGEZwnkM2FDal54pSLKgLY9ccTGOBL7Hz5YcZ+vMvzntjxcisE004H7RBQA/CYDPRIl/ng53
8bvbuuTA9DDyjlhHV0P+9OeesHoHP283oWd40jy/wUMYY6PsDySze0VsoUL2D/kj+WvxEFxNfO8Y
euE9f83C86WlEgAurk/D/D2klIcKZnmyJbpH/z53kwwQNtP7F8fbfOpOcEdpoeES/ctsDPMYiVZu
Sx0p+xzYOHRMMMGVRFNRuadcCqYI4gEjTgDzfLnnXp76mENGQwfG8YJTg7Qs/39M6cJBKynj+hxd
VzCo3JoQRVgJfvjsDOihb4vLIum8tEweaoxt2cOMgm//1VWlJIXC0LRumGpw3KZFIihWyo5Y9+KQ
Q0NgyqWPLiN+wZiylZ1XxGxxGrQh4bSARDqinncc+hdkLbkxAiFW01YUswUqvNaWqhfA1Bvc8Ah+
EmucmvPUVp7tCx44hPQOMX1GjvKpKOIFRBnlGTigOpzHrf77vlZWBZ75DJOWUVa1Kg8QfBMsGHdb
PPSXfGt4/iWstKZuMl+ZNwbHCR58jF423Qo/oLxc3jQkPJQj3EEfB0IRyOppFjdlfMH2gSGpa3fF
dcD6fxj7SrJys9XZHp8Gb/8b0zIDSsaC05bZYLxRdCN7dU6aXjz+UAeD+FdYjAV3zbjrjPHITze7
JqEcsIvcflbtrAG6eQrmj/2Ozj4STR2A9hNNE/SmCJOWoKliwsffimb5GUcqMvvcGFRYb7OoE+dt
7nswHCIaqNPJTxZIuJGR8pzzEv7+lsRPM5SESuCBFZX5LDZ1K1UuP6MWSdDk453q3wIai45fgHh9
B9E6Ly+vIb2os4UvH7sikI8S/ccJt76/TIQAhelABUDUiZGn3CcfILuw46fCFgKP5mE9FWksha2G
H0bgEbXXYrIt43d7qpAyoFzqY2RIuKkK7evDIn6+05tmdROVRHGpFNp5sEWTFApM89bD6985iutN
fo6A5RfLZCfqdSWYBbyoEPY/i40rhfehgfTnH415AIuip0pOitZGcT68Umc3/Zsgs2NBD2KTaAq6
4wybtBEBc1BxhFi7QcTJkpHprF8bqQ03rmNRQyyoDoTmjz7jV0R1OfaesdiZ4YugRRtIdFUbCXzM
sc5Zo4dsiAc5wieTy2cscIxucUGqofwcoZ45GSCrjAyBDZ1te1x70oD+fW4bSXNLGr93rZU28ZpS
omJnEWKVu6GlncKNWNZypfRMVyk0MS6ChJuzuRfLjKQR16tcRLFpXZ/DsFn5PJhszBD7AcJL4fxA
XQE/Dcu28JgXIM+PwUKQiRax7hpDImVbdQ0LaGLYz3VnUQT3p8tVuhuocXnWUuqt8na01Eh2dpQF
1bMLbLAR1AfDipt5Vl+Cjj6bfps7ktrcVhTTDXnbqE2182SiMYCArNXcfxlurYK0v0XbFBbO9d81
xVckdU83BlLuDh/SXh32gZJnV3nRQBPN2vXfq9C8NlWMLSlal+pWoTwj2xJBlfOPpzuToByzufxd
RWYl3M5WSMrnZc27uc7tTWhiRmb0VI9L7nzpKLSiDCElykSUXoCMYWnmrBWlbA665K96rtG/rfA7
p/kBR7F0o2yDbXIFbo2Xnd/kzpmp7g/Kw+omGco5JrWxNxEtG2vzE9EDXbsboIxhZy3NRihoLTOr
FJd4VlUyyIQtiJ/euDT7LrII0Mjb8fOSQNsFBKYSAFe5ScX46EccDwmYXjFMkNzXKUe78AEX7MvQ
uthWURJlYkN2qNdq/tveHQbcCQ5ZdX1B/dqTEWn64NMo3bE4SqYIQ3xmP9Vdp4m9w3n47RBMldQ2
7+mkfpMmUgvQVEp7H3Sz+N/41OtIsz2pbB8PS+g6XN4Icy77Oe/0kyULiXEu5+ZiBfWx/N8cgO29
CF2GON3T67O03dvzEQ0YbJQwdMk799vBvhAKVv49HkxiKCO1RUPkLzb1FXdlRerhMQ5Bu34r1BPU
DKePq61t2a0LlO1qgHz/bf/Bv+zr60Xp2QSpq1AhuAjrCBXMSVpVaVbfCjbIaXR7r46Un0sYhnEm
C5mXLO5x2osIowAQ+PsNCG42q7cT/dvtBsqXWJ0svNwtv/7MHmjintNO4p46a02UxqjoCNylKvzy
BpTbOb+EnMv99XYpENaT0921A1alk0Sj7n2WTtFADSQq2LSiya7gAYwt9o6LPoJHNdHRNDK5BLUM
dnR5l4409P22ISo/rYftYgKIx76/r9u8YUgQiGAyrTt9xl8DZlOhe+OcCvyccmJi9i0mrVg6dTVr
MELq0oKO+h1M4wlF/wweGVlZuO0PJuLtLoSmhHnHE5PQJjmD1yw+gPO5OX5DOSXuNDFXYe7E23Ec
hgmZKHQSFdWVdxJsAK1ZAwX7IGJufKojaqD4rjkMDb2Zw+yedUJLaLL68qja19VElVm4izaXK38q
sMSKA70F0/ygFHDPAf7yrcAi75UxadK9B/l+OW12ZUG6YiGh4tlXvp6Gd8n6bJSf47fmPmRuL5Sg
/cNb/EjyS5BcITLxk0RsTiwwxF+orITrRRhuYylbiY0DabS/iQYqGLXQniApvnwwnXReN1zASpdr
hOCcffpGrNij2wI3b/VT9nVIc1Ygv918QFSDAhjaQ9c7DLA8ccKbour/jaQxZGYbfTVs5vjDKVMb
upX7SEOG8O3FxIAPFgurDZm6vV1CKVmTFlkUTaX+pft0T07/hib4xnyAmp7w2FRdr7NSyZL5dmAJ
/ubHrfqJpHpD1mA0ME0GSwejNGo4d26R82dpYMY+2CiBVLlKFC6k4I5AOyfDf2EwPkaUPQp1VL9H
hlgd15Gk2Ok+MfLFnfL2Z7+bU1HAZRsbIXWfI6ttcK+INe614cABVMBgo2LBMZxXVVBwBSlR7El+
lGbPz4TW0umLGrbfc5ro/AvEEr/j/jIxk1Ou8WsjqaIS50ytRh2yPyHXdrJYpuAtPruQ/VO9q/BD
Cdmnr2cd3hibVIm6zbk8cnoTK/9HCBls/XbQyv8E0RHjL4viYCbJrBMROSUUwmiuCWZGnNk7x7sU
xqEaC+EXuz+cNivnoHi4JRcTnhqzw1ph4HL2lPhPpJ2nwZereCmZqmgfWYVpzYOtWmKsWTXt96aj
axcYLad9TnOb8aaJW1uNjJ0KjV6yzTiisIYu0xJpX6b0wEsW0T/nxcM9ayDyasbZREPWWFc/lB+O
Ddc88jpWcL2h6ch+BCqECsPMJknexActlRJuWbsWUEcU1E13BdPkVU2yfB6z137Nd+g8j9OW2KKy
PBWMuKC96DupWNQSMdsO2UHfZJOCNjXto2xKxE3TqwozKwW5r8J9CDybjJ1T8Q5EOGXU+Qq60IPn
ZAq/JZEcE1s4d+hlFbAby60h5moq0fOMAeeoHpIakDc63qYAsZxYm5KD+TbY86eGhkURpPoPvc2j
H/68kpFOcZEM4Uqz34TEQYqwLYE/48nKABDBXBTLFi76ECc9ZFecZDxkgjd6JsmiXM8YsJ40KzvV
fryqVN9Fu1qMq8eiLBcLU0Ad+/R91+IsWNhueYrWLHxEZoddM4ocroIQnwOCz50xi5VBsXpFjId6
LAkxKlbbO/GvbjmVc1LzbU0qfKePOpsuViGftghZE03T8e7DXc4vREmvaxIfrNbPrM01zSi+mxzy
yJP+j0rOUcpY5AuUGD7In4WxG8yZE8RmeoEI09Xca4Qe9sbV6zzecXPrvcK+4ffYvlgmAj8VY9vM
wcX4nf2pXQMF6vOE7WNHRuqtDmaaTpzimmQI/W8ZmJtiBjEj12F6jTDC/eI2tDNTEICl18yrHk9+
5OgFCpBbhocFMEHmtoh/Tfxoq9aanOUPpc4rQ5MLkFvaGPwlOHwrxDVAE/rfAP+pLTjjv6wNpGyE
nGZG1CIn31rjDi3BnevGQi/1nCnLIPuzwXO0Sta7tKgb7JWxDj4DPSB2OQSl6HrJSMebkElo9Yp4
OsUxp2eivGSKACrZZj9UbE2JPQH/WD9aE5/wh/INIoErjIu//LgS4Zytzy7k/wrJgNk6VcaU3ZYf
rCjnsHBLwHhCG1+tfXCPC365jErgarPSW9csmVq9GBdFmpmIwbw8YB89aCrJ3R0tr44H4Zzdywtd
T6dPl/LpDQfYi4CEEGxD1R2MrG2cLc4zFRKbHoC+YBO+elfGDXd+OFyjGQNpEQ3YqUz+exspsN9S
XQxUxoXyarrupLMIkRicHDgcaU1vRTj+uMhHf0/AF3RtUyzeKTU0xjx86h5krJ1vxitA6wFM0VaN
tsleVPeX0WrbuSm3mFy5heORwvxCaTt1OWkMm6SBZcBDzZH+jV2jV7u4N/uPluqrsdLj7EE4xUE4
dE3cPx9ruVwSahxjpe6Pd0ZOsvljr4jOBnDsdrQv/CuwYSnhO9b0f2Jjizp/mqG7t4IT2r6WevrR
uGIfiVeU2MzTPju6Q0/5gcMXnvmM7Ddibpoljy+twobGjTFy+1+Du+HeESHFLBTbKV4nd8guL3rA
mnM7V89k2+TGst+6aGqlfsEOxrbjji2EiBuYZ/Ekf1E0/hnH8MnC2p+7ju2FigQ3dOtnn8lfAIY1
0u2hx92Q6AIjSlTfH4jDcpzTrahFkwTt3tmb6BqF/GIjB5hTFfqc3Mx6j2nJeus2cOeENFa0Yk6l
gRCQG2f7MCvobBDfy284eXlvBPTLwaz4TRi5D9JwIme4kGSvN3YE3GqEGg1YeZHPfOTS43CiZqYj
czGXRWm9CweAgeJFMeAsUk5/C72peAuh3E7pv/7+kYDKnbR7mDzs76enBZ6Wye6+WC4PgUAli4sp
KTIRqo6M6zGZx0qi0G7oISkc2O6+LuTI1gSufdQ/c/+CvkaKNrldpsCXfs9GBlVDc+Imh0juRsNG
I4J1ZXCfJN0IncUq1ckvUKhEVMJ/IOzaBNDsg26K384ui0Qv6PkENqzpB/x5EKZy2yLAtG9H8rJp
Mn0TP72KZwadMkRK7slphf0bMaXYgRamimLQvOnchSShJ94MCxfte9q7KzIgZgqto05WuZUwa3Xz
loc1rtfIIsFVZIw9YjdeBOq0YWzVZGHBAn2g5HbcTIE5hv8MO90Eop9U+CEfv1mmkD8MAnu2URZ3
OrUQKZQxY4Jiqg6wm9BjjCeMezWgXAlvO6BN4QnQCbXOrUj/Pwcge/IxRlpjvYEC/aPQJKGJyyiy
VtOjfg63vyI4+sewMb6v5SswWjyNOCMcnV6rHnawl2L/HUVOiuaNKKh4qsrp0saz73nmTTMckZhp
UIL7LzadJLUHeHa4HYr32CtO+2LxNRpcNasbczvSk2GV4M0jIRSlFlih1OMPbj66KzrcVzhnhRpD
7coywRtLWmzHS+yQbY7xxuyuAeLxYcDbXT9c41hdR/YvwBvKbLLqMF+oYywYBRDMpYMYZHlILVpw
rK6r5eyf50q/kMKiAoV0BQaFzBUlcHwSeFLrUCtYUOH34JpsKGLoOYrDZSDi6nKYx0LZXcJOeNFN
fswELkbt5ExiJEUuMePeUOARW9tOp7+rptZRHaNR1v3mx88pVNvIXAOQ+Qio70fJNPGu8PNNt38x
/gvLo7xJn3nEhPxmiVh3nMfRxapZH1A9kagOkxADEJ1pkq6qi17afLQKs2cRE05ryoWolQ4oJsro
JDgHJ+9Sj8zgytRsD7eTGURPTwDNXwUcrORyBkM4c7/fsSpsnUJSMURPtS9Aq40exeD72pZlNnXx
iYEq2CshuL4XgZv16Md7LcZq4nWzfJCmiFP/9/xQQCaQWze/3tCjRiZ9gAwNlNoJTeyeDJScZiM8
+l6UVp3FPdyJ9VJSPenFiUGu4LXxjjq1AWtNNSwbqBYklJSdbBaTdL8hAAQ00vJbXAY9lQ4BQAjf
mgTpF3IjlBWNiC1uGrBQq/ebnpHFE/YVEVAB0y1JENX3GMieb/Ks8ZYdoNgAGhBe/TKO2XNWdfEh
lCw1UgQqAILlgdGOHKHqi4rT2kyp0aM7sf7mw8434Pr3LB1jrJ5GVyYKsSkuAc6X9w74+q8MSm6r
b/oYLVd1IYzxs6IHWdbBy0YyTGOgWhTifk4k8Bs5V09o/MuwMf0zroIvbBLocCzjovjnb/NWrUdo
WAsphJe78lHWCwxQ+8OYwZY2y1ysrjWwL6R/s8RqbKAuV3+dqq/cdWhGLBqmHoFT46h+R1nOsWaD
bKMEC3ywSWCqfm7pJ464qWzuuxAivo5O7qgDIcNtvnDvbRrcHPrL/BEA0lOCKBi1MxK0y4waeHnQ
7kyWDfVSeYtitkiUwZbrLAUU3p+vFlhOHema7pv3JtUGtUxKyHFp41WILy+iJkCdhFrXI63JdTYT
2vqy0dLfx2wOr+JzRGaoSka9OAdstjfeUCRglVEZuXcnWe+vHq3mYF9hi5DjITns1wHbfEwd9xcB
oV+sUyWIvE0GuAIYserW0bV6KdjDiOmJIJcb84rKU5XleW1DjRsHKVXxS6nmpe9SG7k81yezSBiI
adaDoAQ3CqurvovqicmbeEQknMSL3LXJC2JLENuVXFsH8131uB+zQ6on8ZtZHfIPIWaH20TKNbs5
ng6rkQE7rxbw5lI9wB9ZDRHQv1p8yz0g4oP7C30+VZJI+gdzXQ2VgM2t6LY5x/0GuQxTv9OomYto
NUnawtc4mWyicZc+ezs5ok+h0yPDjfyEJv3/BzUy8ZZca+dMfFEYXhJXgrEhyGnHA9lxXCOK8sGo
DelS8YNQohJyX+iTRh4cXP6DG8ZXr/INYZTW89B4lLptiKf5aEvHqLeESlj9viN0r4nTxa/JsJRj
JHnRrdX53XQzL/VinBB6BbnI8PlakQbX3cMUiypX2invKJwHJhXXMsoZUBmPnPc+P/QqUea+6uU7
5uq5Y5zxFFtEqeqWdmecgyKfgJDHN99UEksMPpW5dzAH5S7BV5gj6IKPerPxD9V4zHePVYNoluv3
q3CMyddTFdksYL1hUF8p9Cbftgki8fQvaqp+QGlH6YPzq4OGQ80UVGtzDKVGfKpg0CPNIJyTOlh5
uUBj42B6p3gXKY69jdw8R9Em9lcAcBvQvrRrF7M+LQNJAjLWzmfZ9TQAbG9n3njPxPw4kiG9pGQv
6HCOa6i9sAZ/6c9nfnkGD0tIGnQMPiNCos/mNmXx1YsrybQWhAsj/5Ap6alo1YTSmbJKblWwC7LY
L6ebDG39UbjWSXwc9ZTQVWyMkuopLplYJ+QQ6yKt+N9fTgydLjLTBWuEBJDHnWq98TJwKISAYSIB
6HNbgJ2arK42mqRgAm0TVIrB4KLkkFRS98l01HafSYTBH0uNCf3OPnSDRmMYA3Had3hDb6dI5qF7
ZGKMSROIlsPxp3pmcyJrXgf9n5w5zY0DixxfXvF9iDi0fsGOJZXoHjVZ0dkiG7S/uC5uu+Z5sahS
WW4HCzkExJ009uYP/uuoLVJcif8EyBTwdZjUfiLiyucUcrlij0sB8NzU2wjXwsKrXpwHnVh+D2u4
/AyHuoduyxnYeGCBMw6Yith0S10hB6HCjij7f/UeAcNxYq0TRt0Ti3snekett7GUToeRrxqJsEEY
v8j23g3xM+r1NWPYMZn8jdfnV0GP41aE0jSfyDxWekntKBKZ4qRa6kOU3hLz93mMeb2MQpHUAsAN
7jOuBkSsz7NkeTqTVda5gosZLR/bRwjsZs0akAcymCM0SL/jh237JjqXdM6gX+QVLWwscjdVeUcZ
+PaC72U5VJPMAwqdaZUWRv1CyFt1xm40bXwyLwPQ2ysqWL40PzGmGeYH3Y4pCeZ09c8++P7KLm6J
P8HqXMvJQW8Jtt4b1FEaAMZU0wSeudjKzodAv4Yy/limM28cnVKHfZMtVp22yKwcDdhj3WM1mvpe
E8EqEsuJkrwxk2Q09/awdd7wmu2N/c3KUxj1DelP4wFvY0uZvLnGU9FnTsonuuqPZrGwDExM2xAD
udUVXOOQc1Ec//i2TetbTCumjaI5lmfSbqxmZkpOIorwbCyRqps1xyStQXcZ5wK8rlfFiLkSNpJu
+Ui+kwbalCbzhOd6F1TnXT0GXK1iXA8gPuj+9NZrtxoBJvxp490CsbQ/AUgfN0HlAYH6SNcvUccw
LYQtxOHwH1lAym+taMPaaZUIqtV3weqjjNsRXvQbI71z6lP3/V8pphseKnIjycrOYIzEEyNDvVI9
OR5qy8I3yDcnOv1KQ9+3Vu/nGM0MrXYsZbuVYpGemopgQUX6ThLSLr6CscYCwmtqYzZZsbqR8rSD
FW1ovqxabE3agFC/8TNCPfpOrIrrxe6Gzpt60oodlDuh1BhhWcJZnKLMoZOO5yr3QgY3VoPiidI9
+D9h37tPcqqrNS7LLdnF7diCvYhFza4O4RB6oVgzgkp8R28T84KWP5NprrYadPGkeIRkCljTBfGH
LuFjBM+wIKvQQjun0rvuL50WRZH16Akj6QPJ+y3+UguoER+UVpbNaXbphc/vgrOk/UdcKjRPEzHQ
6e42GITuGPRcyYxd19TStv59f8bgMD4cpCVV2MHah/GPCIVWZ9LINSdgfGuyYOygfUzmJdjzUz4P
I9X8nAhoY0hmzspmpclKLiEvOdfuf2nM5Kc26Y6AUQ1S/3YhcoZvzZCl3uHW2MzGB2WYgvXoQJCW
9XMwY6F4caJW4AR/iHmcWSZsrba7YuKiHoSL71I6hLYNvQJ3uy4aKvAKWfEW9lHQAHI8NkdnmlOU
Rp1z79geQD0a4SBFPYdasHP5uGWG+FVMeu97gLMEsz+Cw4l3o/VLvpS1+4Kfh28mIfDKYMM6EJo9
BIkumKaN8UzwswBjVsgzcEJgzY3PoWXJ+DVVurnnZtIXfskWELGKULDx5V4SGhGrErAy68JjhzhQ
5+UzxfJlvFA05CzLryfBXWumEyClZc7dRzHbsP2zJZlTxs/Kjh19QwcSvOC/7qkGo/vugq7OktfX
fpuXppixWLJBWAOH7ihmXzVfybyFDGlO8c0cCESXDwPl1bL3uYryJFAx4vXiBB5+/oYkn3Jn6ufY
hD4MudoF/xQFpJA/cydsyxIJliNzm2C7Rfo4ynJYUVg1OwgQouf669NdqxwElaRrM42igsxkoG2O
cmXTUFiajS4ndcrNXFfwNp4UOMEHefFRWE0YjcN0FwbIANKyx3PK38T0unsrbTLsCC591lAGlqMW
fS28rCiTm3tb0Nz3UaX3EBhChuC57rPc3p+ies9k7cjC1mYgcO4ETNxQCqjbpDHIq+aWJZY3YnFg
1rhdFoOqViJnytXdzV/CTLaHX+gLAU0eAXFZTyI9FHbuJTCFafHpkNPZMc4EH+W8WSF8ouOnMHH6
ecHVUJD7ClMU9M7rY1aUL5pcbvx07OU7VikzL2GVNFc5FRneOV9qWnYdy8o7JaR/9Htj1VHANe1N
6O0uzofkbQkAfrrHcRX6KVY00btxt4Z1eWCCqjkZJB1Nxa030FsbzsV2hi/aWNay1B0dVeP+X8rX
zVx7Jtt+H9sEu+zxXHwHUlOWM/h7MuFtApt3yXjZgLxBdGEGBQ3co0w3LOvdbjcuoeoSfTZGvi8p
tqnBzqC5EMbNuD0z+20XZRwUeuXhcvBB6BTmNsnxn1MFPzwZBC+apcRotiUXdNxD4TSSuvrJAkz6
XcKPlsU411JkqGYkwknSTT7xNLhT1f9FoXPPUkbR6q59XxZ71cjaQ+OAf8/OxPv9osNCMkssSQ6L
ITiKAo2/7a8iNYv/jWFvmqrCdyey272jSWOYV1zHgrkcaW4Q5iak58aOF9iGKCBC5n359Jl9SPFE
l+oIL5mBtOQrUS9IEwd5559C42OPtd//AiCZ7U+GF55/nMu5YxHRCfRNEqVoqXFsnlfPiAjNfmC1
Z4AzcHQfKWPtI/UAWhbmKrsFaHDb9RG+DQXBssqfDaPukaXBvnR7n/MUdk5tItbO1IUZB8Z64pgt
1LmnATMPkpoT2SY9bWyQEjR5J8sE/H+Y7R+fQspdzHlpQDBfh5THDkUkz6/Z/p++8hG3BJyUZhCs
ZEIpKw6E4Um6Io52H0zZWzJu15m6fnNj6zv6l43Vo01LOkONnFDuiFXqF0RfJnxQxXr0e+5K0t5N
BxlYADz/Hv2eOQkNGZ9kE4cpqTkvgthQ+lZzWhlOlgET/x8nxFfitxY340h9/ReTtlNwCuunuhdv
SHSo8nnoGcEEXyVMvgADx2Blho46ACddnaUXw4XE24NYOC8PZB9gUaOQ+lXFZXRUE+y+QT8BD+uH
5M57Sh5oRlf4oDDp2HhbG0JIvd7SW3VsIHL8Q8Z8zBMYEn2QCFs/J6AxF7rjqvkZMPIqYEg1ziKU
QZY0ANKiKkO+xsrv8Leb0eIDtiD34jEFXx7mq9M8/uRdsBQ5QDVfYP8eBhWN/qJH+QrldbW0k42j
j66yDPN3tz39FqLXm5bJqn1Ce6nnUL+TnCWzH4pgk2wGAlO5zTdoFIPhAI6XZlPxOA2IA4Xh4OMX
iZB0AUSMP0vtx/JehTFqr2n9OpCtUmQwbLPXEn4e/0TxejZMLvkaHv0MiBjJXm4Zvzw1sSdoDSr/
43H8A8bpCEyygIgppoRj3u7tAAmVRBIRMM1P0avQoAszIjzXL685cx7ZReG3X8wY7Dg7WarXOfF2
mf60HDcZvNyZ7mZQ4f7mC/7/DDBd34kJcGb3d1CAyW2svmHvsEcnFDbfnSMs8z73EGdTGPRqe6PV
qltrByAQBdfDu/HZ6W33M7EFcdrjLM8V45Lk1kq3t2ZKMTwj5Lv1Ko8SKb0RSVGpMq9pG86yjJ3t
uF0y9BsC8M0WaofHMIdHhPoqYmjS5bilJ4jbvAfUywoNP1jvlXT2/lMCgslvOcltawZKFaU8seyM
XRuNHveD4vZG8bKPOvfaKWWKZ55dpCH5+j90i+I5Veo2n+cf2ilQmeP7+uGz1F7cHb5wmcOjJ5gi
RlmVoKOojsHfmTkaNM8sG5HAGHWXQPI/gMzqmABEROzRhIUdwV9bAyL+JL5l3kGRnGAwH+DoJV3e
r0gd2bLXaM5dmkB1wnCYwev7Tzzv5It3A91S1vdZahZ6R/o+oxwkz2I1XdScafYfQZ0cABrq7gsz
E/MY7vnDiialKVsBNzYD2Oks3l6Q5qg5GAb1Q1cxUTWqcEyUG041lWlvNfXPAwjozmWcBvoLMEuP
L5dbA1cEREstAx8DEGnRcc7yAUVpIx5WqKWjITkWubdOfL2VCJ1Q3CFXuQvwK6eiPApxGaixCU0G
z47+D26kLspjCkC4iWnbqO0HwZ2rHmMZwF6Ti6vHQ1YPdUaFWbvOOxLw/R1K+zPyMEA19x7dxvKM
yffcvv7qKk6eOtA5zismUdni7RG3yoDvp/Jr0uZXF534rGMd6uAXM5zhoGQ8i3tDoCLMgCzCGw/0
aZQ95N1V6U3YMzpOaMfhVG2GF7BkduGncSkYUdXjBF51rqWDLfMN8yrgYMFhy9Q4f6IQJBLXmHb+
uXHY8utd8G9YUbWVC+W8SYJSayXzSXJ+vgMIYTG705KCqt1qGXie+BvrIRauXvvD83mkLGhAVl4Z
xYxBYECJYL6ZkShnSpEX09EDZyg9oTiX1pR1U+OfbE/JymoiNYPPYgduoHrFZ/tqGNDzPzEkEnae
A7+wlEsqn7jgvCCOJLNy66nB/v6PBJNfn8qm0FrXB77VIGjx6i/1x1pAQQ0zkWqUBZRuCTQIG+PQ
mMsUmDZeOKGt8Tn5fl8BmpgvSsnUpYsbyWXCkErliZl8DQOgt4ZAB0YIcxT9T3wVnaNi1YHuyfzg
Ht86wlT6Oq8KazdGksIyPOJ1/+cr1p0ldZ+ifRvrMqZZNgieS9NPEedpcvhWNKAAyG/cMyBn99SE
FNtjOAD6BiGuRqdwSB7MBbiT5QGTB58o2vYp4vIN97GX44BK/jxuOAUz3XTSNG1Mss3O+JzQR367
9Vyf2tHiWo/qnN2H3+WW8Iwue+rXyH5F5Xf+8j73aV/kD+ZapzKq77P1YKEk+qjUs8pr7DI9MjD7
qWDER7BjFmxEIwIzgs1c5l+wi9IOezmv2oseG5CEE5MpBZpAoTOSEpZPGMtoNWcGn7NPldY/TqV6
bqSkUo/LqWQyv+OvdRaJurkW/0phudwaRYWr3wDWvbM6ScpDVCfRlq5fbuBHIpYQ/vKp/pixFh+t
h8qU6RhzegVLvVefRXHG5wnt1EYuxPPe6DMBmwFZjGRb/YK8aXU7F1Tg3l/xn39LBs4ollpItycH
KpEJJDXVsfEuJ5omMWtDcPAqLbLaahoQRqWY4bwO8UBV43RBHk48KmF9R4SkPyuCWq213YXTurME
5YcZpFLduscPYQKlExeQc/GGWBzXzOrAHgo8VtRk0ab5Wgl82mGT29mL7gitt7KCYvAPqHvivlNn
0GWSgJKP9viCQM1FDydXPK82sz+SzxXOPtm47w4laAdAidCXU31jOdOeahKauxvFHkBeQ7HwoDVH
w/TKiGyLpwxh7EWMSbHxCSb2N+N6rUeiokIOjOmBbds1Iowk4LOgSFGCgQaDvuTCi1gfNELrAt94
J1xsMoCaFWyQ24GhML7AW843Vyu3dP3yXvuC3N2sYtLFOIcyg3IDOsX0TdxS4rPmVgJEWUiaEbHp
p0CY/hwLSP+Y5pd439HoLQvN7gPKuj5FgZ2uatV7kEUSAIaQL8dMiLvIhT6f7jjszzcDIaryEr9j
x8fn3WBUFbmHJq16DA7Myct1msCdn2I1Uc7bbVrPKcUZiD5hA2lab6o77JXsUGBGX6eEJIgb19X+
i7BDaqVUylp6KzXtfPNpCbODFdlbpMlvKe4sqKH5JuxLDTAQd9fZeRSKm18HH5JzQZ1nF9R7NzlE
Yn4yqSYebARaiY+1K7QkLLbsMTZHSavsgesuy54q14SH1pb952PnuIdvmJyh9bmGMpINQed5MDYP
twtXLCkMJsImIzyj3ZrtnrohGeefaHgrV2w3UyyZ1BrGje02FoQaoxqOSFmigPlFlKCRYpjc1P/9
ooUfANHSOrtUG2jJl3npdRXfdao81ogJDYpgW3tR72g0YQP86Cxyqt07dYyPsGqDIODD9Ve0l2j8
YPiYoc6uOXyege6lKp27kROVVh/SEKFe9O+ujkOAzjdCxi60ysi2OdMKh0hxpslE/+j+jSOy0DR+
U1id1m531YCX9HIi1cCxWUY4T8MvGrhPctVf0zxV9vF15sfC2/JRQW+XqTZaJJOOQGzHqq1U3unq
A35G1tN8RELsNAQlVrtcFtC+rkT4wR/9TYPd9uoIMc5UaQw2aULlM2qXb8P67W3cKiwpfmwhvc0n
8XGtzJUqIvrXDD97ketrEEa+IIU/oZlIB+0Z0wHwPHneooZT/0Lqx6hpSx2al9Jn61s2cYokT1bD
XGI9WG2JEoF50EIXsTUazfeswopFEKgapvvosGqigJkBzzP2dmKTz+Yf0Jse49wKiqaKIEyrFHEY
hocD0zItd+YnbqvIQ7h9HC3txkImabsIB77J8i/3aJv7S8GNk0Be1lu3PPOeyuKODjY0Q9yDESol
eGBZsS36CpqiraX819zTY2i8wZQqulgQF4nXlWVBumnqGxU/NX8gBKQsCXP3fBNL7698B88Nlc0e
IOYi7MkNDLUwJYLwI1WvkrjfotNjG0zpu4meQMBnhoyHbN/CMIIyjk1cN9e2BsxMA5cpvwn2CNc2
BQSzsU/IQw8qksScUu/xOj0s+cZ1mHdH+NNnX/rL5NZF6T/tkoawdeQaNE6daK5HXFE7pCJ+nk5d
6uQh0DwMrFsxyqmsj4IghslsXOsQls9lvLnTRinbBn6kgdEeN7WxY+zJ+6SXNzI/cOezYVI8tuTV
gzzQqLBL8tfqmlWWSHOjfNXNiSImGctrNNoE0rrEZ09WqIrvAClVleLEcm+Oecz+4+fYFA8wA/Qn
eBMcDBsdmxZYIPjc+KIdpwK6riiLUVadk8SjxVXrU4p6ftaSRbfDUIlhomtey6PvmNRP/d5Q4cyC
3sCHWn25YfpyZDwwNsJO7imXxOXpAjACuCv+vmH25Z6/Uv6Qs8AqSoHuGPvSPdvk7cFXWAMgDnKM
aUfYsWYHhzaCcShei7YGlmIPhsmIh29iuUjjdYiNjgH4xsqDSjymiSldDZXWKnYJQHmfWubPQjxv
DJ1cJ4WK19IcyDk14Ot0THT1mMuFnVWum5qoWzHwgiHgJVAnfI3ms9OeZExZ2OjO/GvDeFLaQGr/
IUuTLb1KC1dhDSxcHzsCdhH1fRbXLdklHp+YtQid1BwOzkLQG9Iya6d17jN0m3Q1LhynJXQg2a0m
Q3HJoYOYuIEESYUrisDL1horW8TuF3MMVo9KrRRAHsWBc3IU/RCpKChwEKy6jPOtAw/RibLq7O4E
MtHbpYORWBccwc7aNpd4l7fc0X0kbY4ZzRHpXQ9elJfXSs/8JoOJEiVRMllFKmXwXkGW7BW9jyom
AREHZA2R1+jLK8NZ0V9fOu20L9B/vtYNUiKopctVLDelr9gs7Pm03SseJiSZ+paklQV0W9znqvgN
ImsXQC2mVNcYSqKqVvXNWOUTTlIIWzCizATjVNs3OwI2PVcWjuDaPL3qC3qYhjMEuqZfbNE49c/b
RySBoZNAt3mFvXR0S+By1d6EAc4YuX+UYG+QvDKLEHTZBjjIxW7F1n+TOnSIAlUS8zuRNnU63HJO
8W8C0qmtC/we2UX88hjY+ZVLpYl/Z2EnMlaWHE2jaZuehdDEvyINRrEAKqgrMhvdD+IzB1dMaTXL
w9A3TZdVZPGp/NrJXTVre+VortlJ1ys/dhpaPKJvNgZR84T3OK57EWJKfAKGOwcmDg+gX7LmwDIw
B6IBFcnT2PaHlMos/AYpeRhBOxuyaNry8ITaz8GRxnKTkg0LS/WIQSwhJy1VnTbyh6VlsrR/JSza
vTNVK34yOl1mq2zerxpKqyem4UUc2YJN0wS6/Dh6GpYUOjt0K4/rk3E2eX5IyGUuuo+zHqIEWrmk
5TBSEDWX9WlbU6Fu+Nlr0rVLEgd/VfUC09poqMmZaFo/URM4mdJEWuIZzJfXZqLhVQHsZgzvCTlT
g36LeUye/r4G6qgly0x/1vQVagq9kljTL1kqzabX0I/AIIln2INDPkDwunmGTOzLzS6NslkoqctY
v2csftiJsJUlzFz/4Sm/o/X+kl6JgE4KxhOx//FA5UC3lR6LqdsAgDjMGL2bd7ytrCDDIwcWs2Vu
sQMzOCmLdsAscfPtdFOPAOX5TWCxDlkhwc1QVJJofT4kwTXxHlWK+JQDJFgQx2ml3hb38r9g6iF7
OcSKzmkUyyqi84Fj7q8N6wsvaO2XgOVzGFkpPzBDNOw2LPkj25ZEAVgLvXAI40GPUgvsrJPLYzR8
mcyzr4YfXSVHei7WJ+jLw29w1z1tu5nnED8jJItjzrvxK7GNTf7f2AQz+vYm1VcDZHYtFqzRJY+w
vHsKIqdmHPIuQOn0hAbM7ltvrM7yo6okWRxBJD9M8mQt5yal9+Cy4kURlrEvZIr1BQ7o4/BnQ5U6
A5bh6llTkkyXsD95ra4k1pxRFStNETICj1O+3GYDHSJ8wRiHemd4zHNMe8E/CqgL8uz06rSct/k4
VhUaoGMLmkyPYQxdVQuLU9OGD1pyxgiWCkHdEkr4UPB+xJ3UiSclCDG8iKd1Ic94Kn6YWATZCU64
yO44N5Qntg24PjnJnTN2iAiA8UNTXA4PPb65AbSyjaR4bxoBvu4xgbO7Vp4x+z+vlIILDtM2Gy+7
2Haj4JEbaTGAmA1YatgUgaoNu5oZT4QloUiK73bn6MVNdA4f0oiuJFKSWDMYY6c4FBcL+gmS5JpO
KVBEGlON+EOItpzg/ydHtoCGulA2FfIABhJ72xVDAodmPsDtN04WXORj0N3Ax6F0BlpAjC4ukr4G
PsjYkCspMJmR3LMw0bO6YboTgZpZ16T1hgKl6PvtzjF+A/PAWJQKOI7jUFlPkYVQIU7UrLbForBv
OcV1VM6Tq9zDqmnTJr8djrwN1zqgkij74YMHpRGnMhhqvdqaD7rDwNPiIR8+7MhNUVgfbuMxMhBn
RWbv1yhiuroVGwnp5oEoWKYi/uMY4XGz5AEb3sTH7eT8WfZdiMpsf91+tRlKO7yZyH9EuSp3SqJr
AD7smMVqWfXI4yk2yyOTHlvMU6LZlJCmeKJXiVLfeXYtCr6dNXHFaHPkfNtexleiINXtfztZ0jET
HmYS7yoaL4zuQly4Gc2UMmOhefZ/o3A6dBXn6LM8f7v5wi+yP8AfrRrVNVRBz3fzOFm2kmS4Sc4t
9ci6DPeT20cryTVAIUT+ieaaCKNaeF4LH//3WR7k8Ba6XVeomWLKy9jlTkcnkgF8NAovDBBbfGkB
1u8Iim8kvN/6jS2Vj86MmVuTMs/oHzKVAB2eg8kt8vEPNZjRmiSveJGZ5691ZLpLAYlxQIfLBnlR
4snpWHZMWPP4SVLPMuvqULK6p8gNSMswbXVNMHyb88xPjfzXdSZd88kOBX8pYpX+hsoOO6SZE00O
fLr1lOqqOEZA3lFUJxpimUK1984Yuf4Z5TZVg42gUoU/a6V+44jMunBiA2MQE4dQoGHyt+jlfYN0
KHyCP/sV8kyvHSYMcdbJEl7YmZ2FDA4eUaU2SR8tdtaZbez8zWWMOwjU5du+Zevcpyfoytih6zBg
NWy2yhnRGyU5KLDWvkmlt0crnGIfGXvr4Es6EhAu9tTGEtJyhw89GOoGedxVPOrYqAfunyGtXtst
bNDCAVtUky3SSwbZkozEAAFgbKn1Uft93ie8kcOjUZVlEio/6pWvWDLiStJVpqOqNURYd/XOqpHI
RwJnVFpGEIg2r6B6WkABU2pGiLNC3IlGg4J7iZky+gqWBLC7t/3kE1iVtlMr5fmXvRScqa60DyE7
wc1buN6hf9R+BdrrlJ/VjtHuA4Y18xegW+6KFnrEVNqJJFrMqo9XSmk2QkCQUM1vEBjIFnxesIMD
j/4nSh4ZIe3ukCJuUaKPzqHMEb/6Q9oEP7si6LfR6LsFWkPTCtBp/4kn0Tv61sNOfht3E3w9a5Tg
KFB6szg7KGJjr9nLDhT6vKWs0xGCYFYUx233Z2R+X+/nUBnJTOo86fQJGH1EJ4SWekrcqmrrffRO
0RGEE/Wr3xLGiRmlfFLcSbZsJ8rmFsN8CQnDaO/RpXH/xE+jpn3opWJa3dwCC1hVa+nDi8kB6mNM
zKrtOTiyV+hi96HUBu7KiIEJi+RcMy5CnxNW2sAeCQ/Tp2xonA9/9kC+uaVrNjJFF+P6sAXu/itE
K96JrSqCe2lSjDdv+DVxi/KOCWjex+uKVsZ4y/MlJxiHaxHx0kvEFX0pBhbedOtQji/bGLvCgD0O
r9XvFPj+jE2FSj1xl4QEZ+m3ARtDiHMUp1NW0i8DT+9kk6wJUqcr9Pm/BxXQOmpo62jDBAWdgS23
v++8UpaRqzeyXHNJlx/GLfQu9Mm03V4+PPUTG345zv/JHML8n5JGP8JkKbQXFmZrU5cNsXcv0JVA
U+bXebe/ssEUD72D0Jk62Al16IAhkOiSijEw3jP5+kETbPWlG5MvDjpXGEtXWwGWsYd3vGLbw/Yk
DSIybbffejNvjAxH/s5l6j54jbN0tTxwIQBKeHSPCcojRBd4CC7jdrwYD5OhmpXgSZdxSL4tcqzF
JJHBSvl/1+swF6QiKhd6MozIYbkFDJILEcA89GTQ4p5Dd3PhKMd6TqtzBYmxpjC0vlQw3OSYsu6W
42h0c8sb8uqUrq/ibgLfgQR5SB0sVLd3DRai0i/Q1Cry4jQa3kWX2fJK4n8z+uoW5IsTsrwAzr0x
d2pfe1ti1InZFtugCN0od+Hzz94aXME+u16IjRezY/NY1tlmNJIdsfF8p7Y7yUER3ghMtJNCF92v
+84VNeGpkWO691SE3QKYrxIPwg2qqfwNZsbwQr4mPs1zofBhlYmmMuO0TSLbPZGOh9FKV2epKFgD
YC1KK3oUNUg1agYOr/c+E4HSTbDgu0TpwiFzSbGxBmjLFIqsxn+pdy/wgkxe2Zo9hO7vT9HZQHN/
WL+vt9tQBDQw0KOw67PTmVPRUAbQS8leoGcyYSgYBHqUUTE+PDeIeP/8v2Br5pE98LQd2hrnRWRu
S0RMCdgZmDERD6stgL1hfhZI1LjrSXdvAks2mIYRbdqn0m1TWNfcqR7BVYEkxELrPMi8ZldUAIws
/EX4vEp8Wp1X3MY11UTcLuuzqnsq1nDfUfCpltK8E2Bx1zmUvIOjygqxkXqu5yH2Z1NyRpY1gTQl
O2aPRg+pJtMGx98jOc2Uyn3XfnhZb5k/UmyPAtyMwA4NusY4QeRXIFYa0qR11sQ1SAMfJ79t8hlt
dobW/govHvBC/RqdXHLDqWgCseekIIlN+g+pT69fNXjHMCDCs1euImMyXbd4F6nP2aUFcmuUjpHS
Q3exYoVXWoecyrLKPEryGmyZJUPclRSkQY454zH266NzFQzhoNXxx4fN/cSExBlQBAKxFqxW9dfa
h/6FPN6fc+2en2BKP0vhOVs8ipYQWyMArcSglKDtm3qKqKRO36cJgRo0xS/Y/1dLaGEdESwfor9Q
dHvioQGQm7iy3QhnI2vRqF968s6uUp/Ph5W9XuceVgtFKMdhLaONv3sB8oOZonpBxKbyQDqm4eS1
qMVGKSQ3bLk/rTUHW0Ertl5mmPfabLTn+c0acO/P071Vpv/CzBGbmrpldUfRiU0YvNPbDbVqWjHM
izeajMsBtEMpOrJnIKmPaVpUYn3PVOHlNIA27ZIjwFJxJ/a0upv2UwUCm2maoQTDL71vCKrycrVz
zOKtjRVXGlshLsai82Uh2/wekeWWWLtesDvFIQJwGbu6f2H7CFQWNcnwQFkrLif12s0Q0nvjJGkM
dGPQCdKBl+DYGbB6Z/n44Gb+Yx6zHRahh0WLCbvfkXYaZSoBmkgBaYYbPqgjNOuGUl+BofsyIj2Y
MaL0om0SrHgv7hqONX4FY3KhLXEdxtlVnpfZ/PCYuaWfXDYnpCusOdo/P2gzNysaotLRnvbk/tuq
go7IcTcSnRHFF0MCS5dNGYkZG2KT8eKYd2gKHVqoukfLi0ZIIv8RtJ5Tv5KIGSypmwQqberjnnYU
4sxn3uUz86j+YB+Mue5Y96v2UmRdtO8iSEz+hgDeEkeuJl6EBrSTFpXS99/o43mx8BCl++g5Mp+9
q13jH7JqJn1C1IKnf4/b05Tv/vM4xpYveOKXWdlKSWTz0tw0nTVp5dQcGeRZ50I8ZlYxoVRD9fz0
YHPUtn3XdwnbXY8HT19+fj92s5MntT+0sAlekldgWsKKtxnA/2R1X9hFUKecFN9B8EE4nn+6qGJk
PjBlMhH05J7o4X84zOw/tK2EuadnlyjivIV+CHbeEvUeRAMniU7FvYYg4rx0jAw6yHjszyLqivrI
aBHZsomjQ8/ObUfGV+YHJnwNArG+xY7NCQ3nuRA4hXCNW7eBYROgzvU95HN0c5Ov8zDSyFbdOiE/
+m/GUKVurVDH83oqcAaycA1Z7iIlNH5cJyeTvRZGQI12PvuC6T4naSU90KEKu5klk4PwUSaEDHF0
mbhWxdeG5mQ6TWSMPZSeizRQjJ5bUua1eLxrzHad6LRMUbyLYK3NxyDNimMhLA9EWm4fbwHXfcmY
LrzFS2xOStvXONUc4rrSZ4nl4z7b7FDNjnLZV27pkB4neshh4/E9XFbtP5blswPQwo9b6SHCQBnH
WRJAO3PoX9WHJfeq+jSzRLWMf/TY/fgRTKsWsXcJVCYv0CJ/k+xxulBncRcvcBJwSG+hlH8mrjfK
LBfihrw+qTKKszwf5rBTbx5Rlqq6ICXoHz6WeRGEOGCZHERAjvxnvpMIivVss8Q/I8Nhdea3IS8h
q+qpFNNA/JoOmZ8TUV+99JSYHgSYOIVwqJv7ApqhR+DYDa+uN1FWkLR6x3xpzyA6RlifjIXWH8qo
zxlDO71BRHDupYolQpYMTwMg3iKuz659BvOCz+PMqlI71jaCKQ2pTzjLsrWC4drZ/fY/g5hMnoZE
L3acgxWwYRZcP/naTsXcNzgA4yknMhGrClKDmSoXijCm/OMwQTi2HyJVcWigJ3EOWNuXxOuGfKi6
BamzHwenq1sIkgD/ay9MBVy0RjOvnoNJjGwHFPpRjjbLbjhVmkbFGrOI32WY2wYjogGR9xnosn5L
rH6uSkAWSLmPHEH5BRfQPUH389uSCst1SwFMB4tXaeUj+fqmlJxbuUiGne8G7tOTALHHRJb9EL5G
APolYraKLe2eAAQAhlAE05ILfEY0hqqJFb984Z1wel2jeh8Bp5X1FKz3Vs3x0dRSChV22f5CalXb
pSpxD1fLuKmgid0RWmph0Jgr9fRWSew1mFOFNiUb3Q0IKjIYCzx2xJm703PAKWAwHWoG519xe7+2
TYHgS3oQrEAvVLZOw1/Uub2rkjp/KAMaJSOj8jn8rs2lpeSeFF81PuUezUvJPfhdYxr4sFWc8m6H
iUT5wGVQp8Gv3ZY+vmE4Hwt2UJAOfMCI7+bOAahhh+P0R/8XgkThX70WdZgJfrg+WYIpTE23A63Q
smRmLtndgy6EldPMgR+Enmhy44aOnSkEfaL6oWsrQAKu0vNeO7uuH5p104UsrSbMRxF6HogUjzTw
BkzJPjU9TzlBpppI7VetRLZ1WE4qNBaHnazW7B8xDySPabmZ+cl7HlOqIcqTxKlzIB551IOkJQsE
MmJOkoRWJ/gj75WBCf0OI3ssfxVwNJJQ6SpNutFqY7m0POarzQMmWg+fp8Ekk6MZsvJVPj1PItIB
Q52P9oFsF96hxkMspVMiPC4Uy5ZWsjRBF4xqm8ZYq+xNz4sQmfyBoyTbWNRxYtXO1sX9EaHqP/Kl
83ettJ0TfYR9v/3ylNPnWV6crcRLjqVr84Zzrq65eu68R2xIANBmEYgGN8k0rybw4+3ecLJdA+6e
dpP4nfXDmTuqSEG/H/s/gN5eJTvZhdxoiOuCd2yHrC0rIzA7km43I7ydqjfz0YY8/sUP74ygQ2Tf
hKjTWkFi7ORJrBd1jLB4P3x3eXdIDaXdll9eR9FwovI6gHkiHtrpu6SpjyypKqOrbZjKEPiyosd0
5vLvQ2BgsWkq7/o/2cveje13k28+PO3drjxC4zS9LvyeBQWudSS9da/W9U7PnwvzQHuGRvAjhWeU
NmUmctIxbAvzuR+6UzcbcHLrxSD4l9JdTCLjkD4BSiGEw2TNPMsuXYFS/R+6UIYEncZu/ee90nDF
Hd4ZNeWPBKXa4jG0NdTz72+fsqF1QhWsX/a8zMVECPedZV+o7doUJKLmHKwxZvEzvPJoNs165AdR
zK/10FVo6r2izpqobOOco+eYz4MdMUeGsWNWyj2tULSbZ+ndhhQ4A5o+DB6LLpRvO/VhneciTF2x
a193TEq2xqm/P0I46iqgiZcna5on3ZnqqiZw/A8bl5HITtLrVkm8XFL9K+ZFDotVxZuLX21B3V8J
wHa8EWAjdHRjC6rKo02AD8nBz0vgNokQ56ayR6A6NB5pt6A4VjB8LBASZnP+L7s6o849R8pGNg3s
Gx1p9hWmt4i/95elzivbYnpkpKxHm8CHfQX/6DBkyqifSIb01xQRLcVlzS+4wjNG3/TEpst0932i
hcI15mBGAJGgVv4zrRdspnfV+TdegeM3wtABnZuw510BRU1SGH99AdHpS37iWk+fLm7E28IXn8Xv
HQDjDLcQLyTdLKJ92gHcMkyQJ1I0DD6I0CBRxWcqowEOPiXGEBFlrs0urKtPNQRLEe5/81xX05cM
IqK7OSLNcvEokwwL6Pdouxd0hBhwywIn6/05PL+GtwBnJPqwgdjSCqm0o92NaphYnSY0fcDjPo9d
WrPGaKMrKxgk+cyw2qstPNzUp7eYphaOlZLQqKclm13V3PvliReEC+2QqzBE0EP+kO51uBeZG31x
22oxtyboasB9dZmph6RLnOxfV7M2QDGjHdCY3Du43XOydYOPWRH93bUDASqkprIK/sOlw1dpLzep
59QGmmloCSG3F4goTWEaMfr37xdDucuGeu6NX7oBq77WkfKgPHqXZS9DFy+wBJ6mY1mONLwB2Lj8
Kgustg+ZxaKnAEfEf04kU1ltsWnAGpPWNtBIOterswtZT6ZTg/5Dbe34RYWfanIIDzBD9QB1MDbx
l4Uj9nzd+xuVkJd0VvsmatZZMn1M3e6mbcPs4bDA9t1JzyIbkppcUSOs1A+sYNRC2Teit0cKwM1z
jSChMgckVuQLpsdUnTLtu0KKqaA+X4mAvxCuoQO4sXEjXoLsVbvST6YdRv0ctvc9pnWbd7qJfhEy
jRi/b430nqJFKTAfY/T6LMdIbKzZGdxliht9h5MK361bIJBv48PkZRE7XPbI1IUBeWJPxKG2NfY3
Zu91EaaQmSqcPakw+Oph2pRnGH8zjVbT9QBWhQ6B4agUcGG1oV5+N9h4fEyIX1TF8x56QakP4UJO
6Mfeme9u+ivvUcgAX5Hidudm8RphZzOegTsc2jDmjWVCvkUTd2bIsGPK3hWumtbeg7A74Uf+c9IH
72NYOPm6+B91elqk3A3VVGRu7CLtSVdzjHpk7KDLZ0eMc6nivFCBTnzle6hEZaOpEEURZ7S+Bs9I
SL7Fy+a/6AdJbQdwhMv0M2QbBh2XFwdTDpfvZbYyJeaDYRRfSNFi5RE439urcVG8OqhpZU5HFRHK
39LxZKI2DtnRCvs/3qGcMwqlFV4hWELcyyaouzewCOYihD8iPgsH2SRd6Xrox5hRcrDV9UktOTer
l8lMmD5OAksTyZPM9bu2fkm88vHK7/4HofDtrb8mhUllMF1J2gLTNPpeO4NVDmami6Wi/k3yupGJ
uDqL20nCSxtE2DH0LdRKBNCDbDj9md/yaGavVqMgtR/Lhclr3LSlfOn8IiAaZQh+tA5SaYy+2iKm
rzz83bXtJEfBfiNa4Cgd8tvxWVvvJX6dbgGLDb9b+Sx72x8b1nWZKEsZRBaB0YznhVmDJ9HRRtwT
xDQmFiV5nCdTDu8sCVDFFouj81URamIOzxCdSeuDovkiOOzvX1XDZhXTt2wpsufVmab4YyQu4H28
/j9BuupDNJrTgUH08+aE/eUzU0UBf7M2WP93OfdNBlYhd4wszTZ4jtyHtqcTipSfQQeB2dPzu7DM
cUqLOf9z5Gg3nBAro75XO5T8Jd9ZHIjx5WG4ZMMwYdF/9EXpkFJDWqrv0P7b3fz/oAGxtOfztEtg
LLRLoS1olsN8tpPoD/CFmAGXmIxgKxf+yYeyZgYgIptRB6aY5162Yz0DjBXQH4jXhjjowr8wP31J
7uT2t/1rWEr6Y8LjtVl4XTges+yAnpAf1SxFe4PwfGwmszbu5nnhOC+xijtHBy8LAfxC70P4x9cd
iv8uDtpVt7ARjMa2tgOUjgwgrPBvPAYixIEZMJIcbOkyZZr1rrpdxnGcXW5bHCpW7kpRGD+DppRI
Lhpc6370DMvuBR4Hbav/rlX88TmKHWZfgSon2atY0GPW3pyyuWSs2ZqZBLFRwCm1fB9/AXoIsW0n
3ciQMIUFLZ4bhuP45b9fjYAterPw4ETk9FH0WT95s5g2CXD6trFwIUEbpmWNwIZihMTAXuv757Hf
mkWfPxM+dSsyz+dyrrOWfP2bJl0CQRjzxpabRzN7sWLIBQG65QURHPFk7JrzRQ6Gak4n3R5bMiPI
zET5z+euttjcTgahv5J4GBqsxpas09eEpqIByAd5XVvga79/qSlm+TJ9sdkvwe+zgQTVO03JpvY/
QrITA1Rcxi2Cx0DJE0+oyb1ZNx4IKDWuEXSPpvl4N9doy5v9vkHPgk3qtTN8kAGGUXp/ibl5gRuL
xiPxEDhIU5wEwAmJF+fEryLDS42oGWOZj3Yj5Si/KvZe19j6TZwb3Td6P3SftpcGiygitrxdfeIq
8BvWEiGcYvSEKkhsK/h2QlZcxEj9I7B302slQH0THrSrUNwB1PEO2AUU8B7lnuvEBOfcuBNi/zMp
YomaWjKPgourTrKpvs78phBV9WL/6djwIv+oL/7SDjJ1o9LGXN8J+yil2d09x34YFa/WvU8iYuuE
jmYWPv3iB3Fa/8rIbJi8SS9c/pPj6EMlLXqVgw7r313XjvC3UeaKd5d/P4yPJkVQgOQTpMbtpdl9
oHnu0Dlfe1HK0dNNpZUxEfxPvyINsmMZJeFx0XoHVJvfGmoq3fRXetATTFjWtP9HS7pugGUK0DfN
1c5VtcPNY7lsrpOKLj6HCBf5Oqgh+3naCuEmiqwoKAYckYNJhnQDAjK/AVDg6Xw6a4gGI1ASaWDy
+zf9Bz6dU2fwHHI0fQemM7Mj81RqDuWZmff4Ds/nAB2nY1xbm/L1/Z7hBQNPXT5BMCLYJF6UwXRa
MvS5GRrNRZaxWC56yrTdUmmHg7Z5KZmRvoCOagKdBKXFQyu5wDwSWVSQXfrSZyCBm8VI/MS+vgrt
ASQQvN+2rQJPWCyWnXPPD7pD6LDDfzkvg/44dJKkzd4OtbwWjVoyJQXU8Vd0ZszHRzslyYXmULIR
2iWKRU40AQNTWDgGfqM0jbPBx4dV8rkD4jlhsavnQTvyuxjKcphRKzyo0xVCjf6FBw97T+k1QvGK
ZW4QnVr+pnre4bka5IjpCcphnxlX+knY303gi/eJtqgmRzunNvaza/5tR794aHuQWgXPzWMYpqxO
TwHnXpZBuhQ91Mkpd3pLaxSkC9OuDHmvmnNo0HFUqmtEGnLP8e5f1MpFk6y++uHq8rDLT4eYgWAs
ROwd5JDer5WqeC/KPBYWAbc1uoBqu40BRWiHpWJph5EtDGdOr080Zv2LT2Pn7KElakgc/Qdflq+k
Xh97bQIjS4e5pUHH7UeyZ92Qr6LkXOj3xHPPS1CfPWNizBN5jSJKqP5/aFX86b4hHIOVEBdM7cvC
kciNtFORBrcFzqEj4drP7YvmYuRcxX/haAB2lCEF6P8IONYKHgXxn65qX6FqEXRr7FQ6whbbHcUN
hqQPmQcjDfeKFhkurqNwvajgkMiBGsrWKKpJMVN0D6D4vRAUZ8ZfdguSAKx84s4726yZK1sDvAwX
itED5H/NoAvp9vpNoS5zXl2WyBEhLqAI0LTZ04Yfb5+NqJWMJXXbxE/yz8DhREatUn91ffWZk1e7
Ma2N9IfWocJytzFZQSa3WpDt8+IskWHVTRQYYvgqPZ40bmGTlWwd7Vorz+cJSq7kc7RaiazahYHG
lbNDKaf5HoJy2G1jyghAwdpipMEfAJVnuKZXXqvaWMFvMTVPVmA503+67FvR0++umeFsM/IAIxAX
71guALzhbaC+6UtxZ2gkpzA4l4eff6FgNDxZHqG7AQnic3iYXsM5Uif8O2Cs66n/lvDVhdnQIoml
2Nbq/0noGYnK00ntPeDBkIim+/xCNiTJPOdayDaloAp7D0DwZATLA+CWbnkIm/kejdfMDOATOkV+
1Tz5XMaSSRE2VDgGee8hOBtxzfejmzu2X/yvXi7myIHu4AtsMMNSwbbqCsoVtpkIu2wYHoaRqSNP
PLO2BA9NQ3fd93yOF0M6hh3ikHZYyvIVuUtqgR6hBd2B4UsZy1sg927e2fGfW+9Cp7Xdtbqb3Za/
qfX9PZTG6j1szcGUTCq2DifEKIHt8ujYt6AjdfJsqRm2+2grjkCBGxyLK0p6hnGFHbXB1jxRprNY
IsApe544j2eeIMvg9PQXCGnCn0EcIE36FxATE2Jfumdlzdtprv8HRvIos2uc7/5d+TSMJN9lq9z5
MC1E+/95gzAbfSfd0z8D5KOIz2KSP5an4exDU9qiNlONj0pl9brDPGhjTCFIzDP7fkeLnrJjhWR6
KiokcTGkviYM0sOIILI7BlB0PnpJ3drOL+ixQU9zD12aVzYm0O5pA4mwJsPnzllcAtnr5CwoXmkt
oAHt3EG5ldEv8tP74kKN7oo7yHUJeFfY4M1r62ocMOEDcKWy53zOeokl9AY7dr5ekmQMKa3bnjR8
cTHvjUtzHbFrPTOTvbaHhrCb8S7Ut2+/BxuMWBJ+D1mbe64/wIUeaFl6Le5wEr6FIWr2p1runODM
LmdL+boP5bFi69suwAJMNjWGFE23hMJ0qzIOB+wKzulhMbBlwHDbev5LKDpWE8vfVr44Z8OcgG7J
szKEpC4bUriPPxv6AwoiLxe1PZHNsTiTDC6iGpvqEZPrqKhpCa8nBNJY9iDzqUXkFEMSS+rMKoWB
5odXH77S7nFef+K2vpXRVqRDa2M5IxevDALw+O1fAqI5EKTq2IkdIuU048Cniv6OYlbVNw3N6ixN
QWnzWOXop1LUhFo8x9vbxP3W8t6fomRb2DSZEPqd1oDBtP6Q6cpnirZclNeQg6oKWcQklXO46ETg
QazeC90rMwz0ckjsb+hZnroQKL9ylDFrIhU1O4IbCfGOsXZiqwg7qiXzhoy3m1wFNjHXFO8PNnyX
TM/eEmjJbxw826QuhPTbvV/7WoZ0ToZvNfJUn407iGPHe7AFj2zMbDtxjAbUpFKy7Fy6DM5Ar/HM
igAh+3b/hNux0mgyUwYobE8XWKp+BcpUPgISpZz6BcIez653La1oIMzdGp22AFOgk6PBDg9TZVga
dnLLutAsuoHqXJA5sB4h2zHAp3FrCe/GVY6pMQZrnAZ+/xw33WonhET29UzcFpplxMaf3VvQpmdX
qYqm00PHg2lteooactTR39/3d2c/y0FSGFcQU6sFtozfoJqfA9Pj05f7y/IHMalZs7rl29pyMAef
5yNx6JCXjkmD2ZROWeHsxj2S4OCdCL1bC4NU5m3OPnRkVYftP2AqRD4cC1KQqZ8P9Dfu7BUYlC80
3GTFbMxHlypbXWPYSNVADFq63fOmbKkC022mAuYK8voJ4kGtHT3tViIg8X8vofIyWisUytuhj9sS
w8eernWE5gg1eZeoRuIKAEtgVt9QzvpGhHxiPKrTfAMNioVX9LHC2wshus1zkJSS2sDpLlHHPMR9
/0QKOGs/smYqJL9SIeM77jzNsG1VjZvj/bdB8edRhWpDGBaDE55UG5455YvTfVpbQwgBzVm0kBmu
EUPe6YsMaF1lwHEnHIRwrQSQ/rt+ihXE7lz7O2BU6NrO/JadRnA8QCrSZ8I4q1ELW8JbPjeV89Mb
sXagLS8i/kdynghqcdrvPS3oSM3fpc89uIE59NcLdVeTvOw1FWvcbyPEIz0hdzABR4BlS5NUW4pz
VqjZAnWAXZmCa4UkFSY+fqZnwITd6ie/Bj6Nb9EchRk8B5DY1N7hF08bBYGuJ7g9botqk49eadr1
hG3/320MiMVpPJFkApL5ZeeJnko0dOuEtZd43tAoqtRm7AKGcrnaQhdOpvBbczKu+MZg+B1Kp1fQ
qlBn9bLw/dHdTJOE8INz0CPd12Z8fun9ho7pZaYsIvxD2mEaEGHlPY+Lh6z+qcVw6eC66qwXaAN2
XfqPm3GWYTIsN1/MBOJReqhv6qad6ThxsfkU+4MeLEDQOMOwQBCL731JqXELUqax/vkS40JDJjIw
mBJRQB2c/kKIOV2VCv+cuOUIIfT+can7Qz7+FncSHqmvbII7JFDBWbf9vAF5abuoIVoDM7Ll6+vY
eZrwRJQKBLprTxVgz3R8dVn0/4atQ+UpfcRaxqjnhfk5kESHr50SA7Uov14EDQo/xPfTJRaxa4uI
awB9BQl5zJUWh8pmyseZdJo1vxR+diZL578Jraskt6CgE6fFu/RzznCcqc0EZNY3vubgg0HportC
jEEJTpBeTkaEPbva9ytMZcznraBIxFy+x5b1hDmA2tUwW9M/ESDWYVsD8WX6pLga55UzDDodR5Zo
aVPwYR+LH6JB2MIQZCUTgo00fbLE4yg/dbbmmFQIR8p/bRnRhX0kA5mnoI8LLKiPBxXY7sH4icWo
n3H1IFEIH9G4Qg4LfAGVwN+wUGkv1aQF+AbssIBXTkBThd93VD+ej/BT54+kdDmRSGccANYDmA2N
MPsfzOg9WTuQWUGBPC5k5vr7i4iMuXcOPbDl55EXeG87xoS8XGCATnpkXr65NyTiqFKHSKLdQyBo
+TFl/IGvCHmtdynneQFRQRlNgaTW7oA+WcPZ/qbLD50IrTrgqjA33XVvrx0N5Vorv0vsgpwcjRFF
TsgBH0PL7xdCWN60OrlKQ2PKimpgIlPoicWvZbc3exJSeeeZ6MIw6QR1MMxBvasMpk3io/17bwv1
vKMhPswCrNzF9GHfYXwCNhj0dzESHviI20p9fq+W9/fHKUi2L+K0QevWIFaiTW3d0G2rgY/U/UF3
vpOHlEeciZ/CMacq7CZg4d6S0+3qW1+KkqsFRk862B57+6br3ZxGQADqAKXMmYBL8UUlc/PRFRaZ
Waq1SYH6RhyBsLa4sv+2tUmZhnSMPXNkDHXDPfXHnCMUezeWQE1UoMxl3DgEUPQhQ0ONeHejr7pV
egQ1zHSXRcoPMFZMmWPfRKopNaARGXrjJ3C/RblF7WpMnXBA1migDo4BRKlPKj/0t86nbNEcCZ+p
NBqh/EN/DQOXmqanO9Nxlb+bFyATAX/jg8B/Uaup/w6A5BN5CHTRE88Hc/AHD0OKzGW0w3Sy/rtp
IRmTgkwIjB64aKUv9N7ENo4mI3agJ6/7Vxp0ARwpSIK/vGVgbwIUt7LzKHmMLjjmtykbpbbNXTXn
5jzc6Mz9RGYwdBrYvQldB1JCmtT+HQcfZBBrFqLZw2UkWJNRwKWZHJmSl0skadW1DnWYJYw3a58J
tGxFK8Sn5npbQR446yNTux6LrIdF39BOB+qlb8OsUMep3jQ+LlRo0PQ/fpCoafm6dxEWTMtZ1h7Z
ts7tSr8CfVpynR8YwamwVsTwhVweV6t8bnJCduULzmwcUbQdq0f5Xdu4P2Tbg4v3/Uxz8zgmtsnP
bHN2RKtqTrdCxjzhVSfbGGrTSY3fi/Huast/p4UnGF8KOMyGxf4zBsatv1tS7aEb572j5naEsKsB
b65jfbOtAaTsCXNJPTsuSkeh8EoftMYTphz9Zo2eJwhkZIibtPA5RchR7jA/WUbEOrntSrI/OFEk
PPOAQXisUORIgJI6ouX6KFZBCw2F+b2KLUKa++vrvC53H40vzT26bZHrL9OdE5sTi1bjTJgwUju9
gCf2JtTaaMo5sEqbX6J1bJoEV2LgauHX14B1QR5XfFW2qpu9VqdjGap3qM2MXl6axt7TCbQCdTyc
w4Yj7TmB0U7Z0FudxGfjOcFJLwYAu6sHNK5RllwoWiIJc//BTZVoSS5kWE62kaBRASxbt6dnunh5
WlXkFRXP3Eh7Rrqz8o0YQno9OYriM4YP+NOuXRmvB3lAuSXOtnnMZxDotGw/uFW+iyyDogkzJbud
t5jp9yw8rxQofMWYFGmbU499RqkxPuwajBZVWnG9Rn6vLDfk17gMe8Aw3U//NBe+PDcpR0grlDFL
B9sDBAPFT148SBvgOC1v3mHfrJgtGTlbBpTPyvYavfHyBqxJKUJbWhRkdmEybS8iz17Hn7BR+2Tw
VJ8S0fWppYWXL9R/0/LwlPmCH7sAIloa6ejv7qlrxBtJveDkiphOyZMGx3lLz4q0hFVAEpw5czY4
F1zcj4Hd6s1KCwxF6uviFNV+03ATZcvpOBai9qp26Lj2x8fZyrrh/xTkVJxA5K5G8hNsdbIl/CH7
rrZ8lDy0t4IN4lVPJR46oErCAhapEHFz/uf5Qf2Rw+EjLfL1VtxU/GUe8E6ynrGTAAbAC2L6YrF1
huayQUZiNCj4d1SCeiwSCm7ZMsnl5AfB6o1uhJqe8lMcx6/XcThSOyJhhFrHoznMyFFwCkIoA45A
GrWWoysGKY1qiysMX0SRk2OtPhgu6MhK9bbPGM0Kvc0c9IzsDB+iwMWEJUHZl88b+u63H9ZaVvlt
JrtMzMmrp5wG0DJtRo0mStESzw8pP8Hj3ujh7X/P4e8zFUqioUgJ9aiMQsfihRe2gk2jnBqbIl0I
1DeU9bfjPApsO4izdFPtOmfHPi/zECvNjKr16Kzg2I7OY/jI0RxxyombJzxegov0a+MXLgdUy1io
im/S8Tcjkv7NjzjpvVkQPb3nZ7+fwWQDeZ+nJqWQAzlseIXsVs6bTCu95f40iTINyA3ePErYqrqR
b15nzX6hfG+3Kkx1yhLYBnqWlY37EayFouz/x+0X0JsZ4kQ7/BVtGWx2dgptuz1hlvoA9U6sbvmM
AupWkwmmeKzhswvN44iZ8J8zdDRnGWXn2VzbknafsGsu4RnVVIemGaFi5/4TrffvJgoK4tyoMJ8j
8wpm/SSXrrLWTea8O/H0Al0cuUmHUrZ0KS8/AvnsWjrQtYNis+fktZXcrQ5aLpBudYASuAmxwPP1
ozRevUSnLZyovudPZBHDR3Y7bAOdAGdVy1GsLuy8VrWNHlaRJXvEBxzppUmXMZeQ9M45nKzrnX0S
3zCR2UdbBtzeoS62jDOMFTsHK+aSJGCPJ0YTHJmUxf+uRe1tzvZlpbvSvlBNaA117SjQhIX0Qwq1
oH1foeFs9/XC9MOdOpU+fPrNwcDIfSFcL9d3jDfgkFyQLRUOut4JFG4ruB4ju1srvACkXX6y5Tjv
dPXKyD5uV8QCZtYhwiDnVaDYXPVyerK6HuD+Z62zNy+J4dtYNlnV9Eaig/LdHXfhZB4e051/1nFI
YgyygssXuq0mtFUD76E9tjcJ3UzaVHwxheCEjEviXu/fV2rbpvE193HZ6m7JrrXIk8md4krqLlE1
Tnhpo8tknAL82r8ZPQI7qddNLLPMjEW+rg7LRXrhVZaSsOLRgVB08jNo3GSdwSsf1SolbMEII7Mi
s6xnWrrhaZzIK7WwEYmipc+yDROMc1ANmbUAb/X9gGm7ONg+LNBkLEc68Wzry2g2rrzvIFg8UrIL
g2kALzywd/35xjogS7Vt7mDDCaAbVmnhDvNkM1I2Mhg0n6Hh74cFmoxKxWOchy5isWfn7YLo3hb7
kOJKsCYoW07LxYsA9XBWkrSenqQAkr6rvSCUrExK7ON0uH1qEBu1k2/2DBPfrw2EwThxrzF1PcSv
UZaoKrSJL/t/fqR8MzUcFPIbWi1q2RpipWExCgI9zxVmzPdsI+dQvE4obCT+hwmMqrpefDUFX7fY
HdMgq2apUcu9U0w8gQ45N9EQGH6y2EPi6pIEP5oWJkb0iOttXmFuJtbsrGhOfgMirhAAsKMxtPEK
2nUbxI+w0MgkaeAS/Jjh5QTA/SgpOA1NFts++FP4AzrH2p7rcZJzP+hqZdVc3RWzKTA7SsnQ0/5b
1F+hKnu4FvEvMfD0LCBbjoI6updc1c9asrpHNEhkRBb4txZqa4p0Vi7Y/ckWsGtjHHn78AXjFqSK
WlejeE2Nj1IPkSQYkU2lf5fyz3CSHLMubSycMXhu/bKc4+JLwjOE/rDCM3Wl/cVFo82hUW7kroz/
t0OLTaHK9GFH2nwJs3wcHQhQl6jLUTSRqHwmzEyA7NDFsDhtKonyup5zC3x5pJ6VkE4J60FAsRoR
5qABGpmUkZ67fPPTt4RFr8f5wXGgCqZVW3hovSu36Bc4UbLCAXUQ1pePtvhVnYXMo1YuKgf4l4j9
Hk6NvanF3Hzo+FkJ6SOpqOh9F8MWtbagbBRhZPG7ouJcwxM4AnrqzbbAFzxDvEgEy6Zc4r/rSVaT
ZPP4gdodFkr4Uew4trBaRqs4qFqp2t/j7VX2ECXDGlY6JvPQWu0e6bvY2SmCio2Zpn5WpoZemnZo
OEGgmx1fATFAXkj/uGh3hpayN244JLyzGKxOpgXfXtiOVEZPnOv374DbRuXPygF6sjEs6lXLH8Ma
+AS06Y092pCSKuMF0dp+/I4dFwh4h9YpEkGNk+FrryF1uXFVkKYeu5Q1fplxr4dqBdLwUTm1r1Fy
jNLtjoycLh8BiNa65hoW/59ILHXw+OtKAesgl6dRwBQHs3jROMQFx3jzR0RZH6qVQaUsB3/THYcT
UJ1VtPsqikwW6DRHhYZimNI4FkboN4c/m7SBkSaf7zJ2gUhgFcy2cl2gDJeWxLhK6n7yvX6slICC
1dhnNtUnMelV4v1J80DDueZHMpUMEJqZkmqtNMMQ6Ow4YUfwLSQl4ouwmW1pNEO5zlTUPzK/gtCK
Nn05hEXl3S9EIKJ+QddoY91z36DzUWOvzUbSG51jcfiCfFUH8X5EFdAvyDhbHOghKUiq+R8Mpgj+
iqH+tcU24tW/7aQz1IRWbo4QVtEpVoItZSb787nznE9ZzNc9vslHBbt+aGoN+RuE7iMR1rc7yxGN
FzZ0LB3BryJ2YTHJMHj9NTOL/FGhgv7yIcGnAcl0K0Hck8bD1p1sZse4ddCgMza7QbjeHgC9qO1N
tFP6HFDGw7v7EyMiTJx3IjoKTfZyX/SFEvchkmZhCRTaga/vXv2zYCoS5+Fyih2UUb02BpOCbcRV
pCTEMtYWJCGP03tOb8oE9GyOvPys5htzpgnthoqHuWL68YGytinZ3Rq3UqWW/tnL7STEyXi7xgHm
SRJQNes0Re0jt+QEnzAgepZeD1RSCIhR5m7Fg+TriW+CjOn7HhDkQDAp9icifgouu6lpgjcSQIVq
CmSlDODehOb9yF7Jmtc8+dbQuWJoHtlN7yGq0HQYnZVJQgQ6T9guitBnsWwSFVxUPoGUU0u49uJb
E4L2SWqXj+58lS2FB6iC/PtHSgjOL+xn22CxUM/7clGYfupm6xzrhZ6h839ydof/GiLuKkoxRCH1
4dNe6zTJxAn0H/KCllLaWCcXQX9sAkLCeswQQCnXBzDvjepEjJk6yE0WhjptsVa0GLM5Bz5zQPGD
WTMe4YxtAJ2A+2wTa1ZFiTfnQYcnHWU2foKTNxkSxSmJes+XgHFo31vWuTGnFqnF1jPxfaoFzCQT
CrBC8Hocro3DplKhqLbNJrc46V3iBbqqliJb7SXr01D+r+8IAOLPitTYe5JM/mXPrtVtS1qYkGb6
fHRI5AqF5scXIuQAXptbe31IkrqxwkC8J4gYstNgNVSl1oIViiJMpuVYYXUM+lyiQmQLnevhV8PQ
IcR08D37EqwO6AZyVdYwcafN8ZeW6SZyBk9xSrwtVPcWTsoXvqKHDWhdybua0Qp7QqCvmQKUychb
hc+F+4WN4Zpug1L7m2TF9P5gVuu82S21Z62B8/qHzTdmfbfWNtdgwS7pIkaB4OfSz+jielFrYkL2
exqSRO2mOXFETuZ0H+7tK6hT093UHxNO7WWnoT7VVe3oeSGq7AoaIpFU0fkhLapI4Ipoa1mPvSdb
a5m6hDQttUVFZUciJ+xsB6vuQprwEOHAj5B50aiowbFli7WSyMXehGiehv/vK2l5+6O8qwjMhZN9
0DDzFEtp8RCfriC1M62lHSfobOAdos5e9Ng//e9tWQPzZz2UxiMF6wQ2ssz6oBxIwP9e7lRRi+Bx
nLxGTgYm0hNKqmBozgTgQxSecdGiTa3hDyDYvwobPfOo/RchnRN4DvtgqfeBaQ0QL5RhAaF3aRBX
mEZqN8IY58fNcXU5ngMJCceI2qJtQb6b85ntP3gbhTM3hDzfnAh5qiM/umNq98ZwrXiJBjIx/rM/
hY1ExATpRWVzom0FxdNEZB6y8/bdHxndW0EJfbPJ1ocw9UprDjT/04c06FA4g2JWORnN1Oh3QDTQ
JDxq7STRa6CV5lp1/NPT7v21FjLm46gNu1vrqo0zmKgQ+/vVWhbs+6pKAk11X5UTW7NbwPqyUui5
NsGrA4Rt79JVvPGWMpcTYFu+RFU/Acbo4yQPYBpIhQNxHTkIPhLUz56bJx3HugHJmxdqNrFHms4X
TMyu5Tq7qHaXjCarPoXo7TQZJOnC3b/lDYF4UEmLiJywCZg31ukCRYZxDun/IMAHqkEg13A8uJHr
QaPDdZa1vYUjowNMp5XfWQSUrgzGqyOnIHC5P6YqLN0T7hwEn6rwZXX0spDVNxBUDjJIOtRR8MQ2
HSYBP5MprMHCLREanGND5jpZX7EJt/1mkiy3P4RIrk2zso0PtJqOIOs3JidYloJh7AI/hd9G0uZi
CceGIn57CVX8IlK6RoEX4EvIHBLEXVKgEojuTaMLFOAv5bPLeVGmw6Pi68hIR/QHzScF1j5RWdm/
nBEmRwRZoxaSUkTXNFnss/NICdEzHHXuKngQX+pCwaeKhHgS116qz8W1TPWjK0GH2oA/5yjZHJIx
VlmiYaJmWjhpCT2BOLnb3HNCIgaE5KyiXOvurpRjgCZXTaOq3o/FTqvHW+X+Wqz307NjDt029f0r
zNOwXb7geH4DrcGo+bGRQ53MQHqxwBLQMrwe3AeRiQnVt7czJ91W2UI/B1HJXY/GvQFUYRYmN+M0
SmGYIs4OEkpui4rllw2w5PqVaG/XivSIW3U9fscYVJjUXG6g8diSRZVY6LaepJrzfGP3uTK0FBBR
/hXtmT6ImoBM7clb6hWue+TaI59VhBcV7YlEvFWeSjt8C18gHlu2KHtww/+HJX7L1RFO78KgtwqY
vOhJLDApBoDOJ48nx1x2kl2s/RQukD815Z4Aw9ESRIYIJQ8RR1qVuNdaFuci57RqsJQ7YbvxA5+n
3wVmR0MpYRR+5AK9dhsEYYEad1JurIcVAmcchAjUxRfSu+j5e4Pkh5JMAPoOAhXUUmHVgfql1orH
3vcWc2E7QHCSy8wQdyzu6W1tOw/Y3s1uqzESAzXyCFfyI+lvxUxXBr0UCuv7UhIav1D4SEBM8eOj
fZHq8vJDZwPuPJuGSXASwAAHt1k+8qxxRw/Qz4NQ42t0ppZMWx6Yx3hSFhuiX1cwnXjztcXMsQyD
9VU/ZJJMI4MppjfM1ROjuMt/NB0EEaGts5QBLJlTScw+erNLKtPDL26zR4CvNCqf3/tQHwVi4Qb8
bVKQbTlW3qbVmyxcXEszrmSaBJvshh4qAs5WJ7KCxmHnXoeoauDMWYQAD92cXoHUid1+As5pRvj6
/TSAqXyVB+1RsiL7rA51a/5urwJitQm6jhKoaWdPsFXw1N/VJJb5Q5XM2qL/+fBfSSFcnIjYJDy8
daSMCcTFGYjDpr0AQNlGK+om36KR7RT70W69CRgiRbMRzmao2qmbftta5gDdYaR0eIN75bK2QgD/
+x/pZPW5IhNc+AwIlxqC7r/bvy5KyrFqrev8g/4kr4t2vf0A8vmsvI4e4QBPw/j6fN/bIQjwWWyV
eVP7bgtNUyhOGVbhCyNq395UUdnnbRtjLF/djty0SUsrwHE7sSTASpm49YL7OvEfZA11H/WUlW9E
7vQrv9hkSnBJ8OUOUoPxJZ0txuPxh8FZ41UJGDPdOGTiNA5V/rxsInro2+2FiqU+DJW1AsEbeiyV
13TtPcsQmgOaOPvqBe7v23rz/53sAOyBA7SdX8xpX6/uH4PDXyqnTQkk0nKVf1B6gTyjHtiiaM/S
jPMb+TEUoLJdh+hM3BsJDFRN2tIUiVIqoP+oxuMvJOtqGntIJ90bw4xij65tNFMTRUkb7vmldsjq
Fr4DmJSHeTLnbiATQH2e8Ypilf2CZWOAp7MTWqnh2+NMBvbr3/wsCdAMjUOIT4RInOAzr0d3aSa2
iT4D1cXECtrQFrcV4Qb5SAEDsA5gYvR7ITjctI/NnrXSyxZBEllm14rzPhP15ndiRaOGlpAa5DXK
OSglZuqvwHLNR2EX+7H27yqYpWbi2/gsm7vJlluVZbq6CiGtm24A8c5EF1nzs+R7YwKOIuZXmCep
JmmfYujLO83k8AktoQX2eu2n5BMiHVxAvx+TBZdIUr3g6egr3uS/9AhxaGC+D6GCmBKQouQHsPk/
PZXJUeRoNhDDrcJVA5L3vxs8HXRWV9gxuFA5zagIX5+m8gGXejKwup993eTqFJ2d0cdzBoSipVWQ
VnyzMjFkl/A8LzNMw5EqA5I5BtMsORSEcM/lUfFGBvWFNpIflcmC/fMx0+2KGqELOL+MbodYYgAC
xXm+tDlouSOQiIVgHrhE2OTOIugcUyzipxGM+CcKaMhuuaDdzTo6ChtWA+ejhlNEreoKokcjV+aD
Vp9qYLR3pz+fBSXnts6gXLGYHxlgoSFUqG5dRpMmlXtwDF7NF/0cZfCV9svyvbUW5MURKiYYaYfM
03MLoYsDbyO3WcIotw2ep5UM28RhfCv0ymWJzMqcKrdwwgvtv+HOaIla9oUayvdQB2SI0kpxPKnp
H+9LXwycS/zU8rZ/AazXU84eE2wqZRF54d9X6dvha1evuHUcdnT6AQwHHKC/KbJLL+W4RL7VXJps
1Fu6/QW1A5vQgLCFxqC19TiY6gQrxfz+4f3/zlvVIjenLE6DvfleR+E9ex4cw38AVMCFrYgk6aXh
dFGwQeST4r/fk//6bdJDjdWAcbl68NQH42bq/GPM2DBVUa+Olygaj4vcGvWzoTfZReixrKS83GpJ
jtMZbpHsiSmCYE9nMVRakJxKC9dpT3X6getdODLQ4j/+jcuQQ8sKgiA/UqJa7jolDxRcpAYA/P6r
CUwW5p51s/jPz88TzCYb96NS8vma/JkSGi4idgmQODq87QuJfufweYYGfXfy8ixAYpBLKB9VhRxR
1CpfeD6DGm/Kmpq8pr3E2Q8nCrNBw4q0kQ1h9xKHoU0xMvThHhCmGnpwpd1LgeRSF5p8N8MsriVE
poYPk7ZOzGdQidrjjrxgRtnIa5l3+nGfmwjUZ1onilAnNstvHdV+/p8WpQJCq5tDr6JMnAuuj9TD
vpA1W7Uz4l5pZnfEJ9sacbzXuO3i75kX+SUX082kBXMX7VfjHveojfs/56OmOa1epMufJxKpKOiJ
pBSqO9B1f9gI1/oPb0LBh1ySFfpzqTZ0kdD0gNf65Xc+oFHk5KUGHWwg847nTf1Iiso0zwRd0351
owiEkwc0w2jJhmSQrzJ/19sOQRgAqE5IeRneKxnBricn3xN4hr+07pH3jHgugBQ0gUda1bum+GYR
pdyB0mcsyQLazpBaFhUFXmTfdtPq7ZsSe6aVphsI2I1oSc11f07WtBzpusvfKLV3ebDx6jhul+pX
RQFC0ne5G1+tie/0XdXz8PqguviYMP4fCQ4RluEWGxVHvTrT9clPJ45BYLgXRhPXv+BqwE2yi5aq
Efa/tGZbuhV3yVPLdCN/2C2RviHLtsByttBqrBd6uh3IVG/f3SMzRS9Ap90Zn2qW31ypvNTvjf41
aJH6Bh9Ki8Tb4sC7iQOcS7JPZ0DBBWOK7zLIBcdxmGlsKzUY+siKRUrLWL8V34tpwrwazhJMnz9l
/Z+GseyIQ5pFw2xzCJYTO8TJliTvfpBPsPRAlAVdMPXOwWUS6Vn+dgDGtKo9BD+RzCdu0iqqz4Nt
iJoRqE6+RpGSi3MzLYuHwsQjb8bShp01+WpNfUdu1260Ow2kgv3uI1u9JbK8vzBKbrvxiPZZOpDk
GnaMenV/X1j4G6vqgzEp5wijKA7WFYlJgaq0QqRL+kI03LRIs1Vlx1WMLVtaBEp0EK+0cAMOo7rk
99ArRBEHVg5Ig6a6GQzXYO4CUHexqcO5mHwmrXL8kozCPlJZoKSi6fEaWXtz11C1V0GqyQeAtRiC
5Id17XsEyhpw7J4hmEYo1kDarHqsSIL3bxpIR3VSO3HqySH4/MPRhfK11UQQMTlHoyDgK6Wr0f8V
+/5HjoDFjEegmnZr9K7PEAbu4zAVzYLD3dVTgqwkg39Ipx3o+FjImnF+ZiSMBLKxNyC/dUNrp3lc
XglSw1DIy+Q0E9XxD87G52Q2cIT7GgHZjdHhiYNa5WnqgTRtREFAppB7pg8XQWQtNxvpbz/U/N3u
Tw9vAbLbn23UNeN3JVGwCQLmjtw773QjSXiiyg3HsHVDcbuzKDZ9xYhFo+LhQ95s9ojOvxIkP6Uk
7CpbYaH36pMTLxdddLX4HfxqVZiJlOPSa+PIGNq4HvWnx5rjdNOJlNHmh3k+MU86uULUrUd/RCep
cyQm5kOuy/JuwsMIOGesd365dWjaMTnuiIB1QmHehg6YC6Vblj7XKe86O12rVJy+Q3TZ+88XtIfF
LHXoiNfzFz1RnnC+//Hnxh+ASyzEveGK131peuQ7ISJad9Wn+PW2p3BkxJ8EhfiOvJ7+WAaFB6Pf
Lstq/BuHuZDqdUGf/ARJi2okhzVur6AkN/GaBecQgNEdZvfA5F5jNuwhoqktfkApHsxtgoJFChZW
6PHIFgWu8MbCFOCdifF4wfkVqee9Nrq9qQayhy9myKqo/L4ROOzz+JVp5P60R0jF1AYpj7kUh+RD
sU4lo+Mt5yiWAr3xMLn39sSOHsFd6gP19JEIUy4Hp9uRm5b897imYjMIUgjwRNBeNPhy6XdUg4BI
3QfRkhdkVkGRcnPOlEmBf4c/d/za3goXjsjUYs4MkqkpmXpXNGYPmhSg/2AIPimf+5TY57uAlBQF
R+7BfpdFoLhgcUcs7AS7JvZRGS0F4nf7z6anRrH/TXhwLpa+SH07XYTPNXuO4Wc1bGISze4O+S+b
chub15RNcl20N6QlS6r1bq5Z0nO91mKDK5rQ//2fqS/dyJZrBHCdH1aCwmeGTLO7F3pFaZu/boAL
D1MRjDrJgXE7rRBlNml+g8BGVd6PudnvTDbwxpOoINaLqQ5VpmgwJZ3lHicsSWFqOCXBtqlXheUC
Vfgb6dEcHST5irUUsbUBl3vPCQrwG43cxLjmFIQCEd09P4g8+kQ5kshBb4LA+NcaHHgzDVFpVECz
G+Cu/X2JpNSDzDB2lBNRgrOE7QLd7jBMfxCxlqoKq9jmuKKwk/SXa+Q7+cyqXPpXkJVTClCCXUSt
xTnyKbA5rfXvYIqMcGXhZQHyr63W76jMzDN1cAeNWD1a0OfBiEIpQwTvBYTyaE/YzYHQnHJfohYy
LBapAWt5igo/qG8PBZq/AHZQf6TvrL099NHRpzotz+ixJ/K8tPGW3jeeF+9pZzj+Ez94OQfNgyLt
Ccm5LxP9gTOowpI4S1aqdSH3ImbZSoI2KVZLCFHBQcTsdjj6Ze250cFsqmq7YzMb/F7i2f9oEH68
JP7dj8AVLTex33u+dNhSoHpVikyxPPn73euj2W75k/iybWe09VVwnwzoEvmOGJLhxA5NgUrLwpTI
kVCQ7XjT523JC2HtTUeZqRD8710xaGQuAVmrISOOY4q/LfjuPllAugAZbAw3bZmXWaylpd2PXYx2
nczUdm0/PXhBcRDK40xfS+HmyV0aXPEAlySZyeTzbKVf6/eb4yEaBoyBqRCLibMg4WwfaaBfOoiW
uLZ62tOrs7nr5ufeg24YU0LqbY+H3KCILG4vhQNRq4nrn8BIGe0wIrKHSAt+l1eEo0xNYpejs3Sp
/IypAItp6zrae11R6hydpTpouYJduy/SDD60RM6Tgb7URw4M1/StlGW8TbNRFRBV1CZPiIARIA+B
0khtd7Nb154HAXOOuHDXzi9WXTdX2Xw35BmMtkqLvnSOKJHKtZBKpZiEFnyRrjr0nUc/QP0+AQBm
0pPAYI0oXAliST4HCps++clwIIipP9ScZcd92VrwFSBkOABw0sy3EaQdn5KxrFeAYcMtJAIxlM40
B9TWiXNfD1emxsu78exWS3YrmL+jHsoRV/jxyJfK1xqMU72Oy0rlWQTpa6vLni+I2eBftlBtT2q/
mXo9U1mmFzpW7yZnDk2z0URdV6zj3XF5BceXzs1j2G7M3D5GVZva60bkn1XrSbvl1rZnXzr9nQgP
WuMbzFNrDW1TlXGoVo1f0XMSE0gZWmvt+WAGgH3M9NCKLCeOAI1rTtASxP6NxT4Q23K0ePxsyp6y
19OSykHwlCTrdmKDYnmOhzffcBRCjQzjNmYr0qyDOLu4f74Lu7OhF2d7Xr051Gv4qutMzdC47+u3
XdjyOU+9PtDE1Xcbvu151wGPGzvcjR9W8+0EuwnyF9kGBIhKgHQ1m5jC3LY8PRNRGrVN/kNXsUy6
gXG/Gxmp/J0WmGaQ3zsCFBwVMoBVZHDimIjsDVQorBsUbQXz1Y0iyxa4Ypg8m7xc5m17jkUSGJHw
0tcxwPtJcnUsJB4pUr+SjxTrTURGkVLCNPNrGS713WbnHZyjKgH3li8wVc1rniszYOdXJwkR9MBF
d07nVta1YVgyGhgOY8Vho3INvvLVGyNV5y77AEAVIAMRvAmYJc4ATdYfuzr/3RUCdP+ycKwxbSBQ
KGAkuhpYPFRoAmzhBY22JdXjVPxuHDoWsJVgbo4A3qNsAtzsjGwC/0uxokOctRd8WWN78mJi6l6q
4N1IUAI3f0DdGBnEJtiyovtZWwy2UExgrPORV0NGoqJpD0kzpYkaDS1n9bYiIGV+F7r6MKXSOg11
2YR8HzbdmZi3KN33WIBmQfdk6mEQfqcQXFNDmLYYwfjLmUArofpxzy8s6poa7Mh/Y2yCFhFkZNw3
pCrTx8VDscpHJM5K8BAPn+p7Y2MCpnH7e7luvl42qy8y+vtWF8iW9PmXiICPmEnTp1qrMFHxqlVu
3cxbSbOq4NbJei0wWZULNV9nHWut8R6aHxp1Tam9qluTieW1I5d1qzCSDkban/jm4m62pyc+yB7N
iY/RGLATPx7tST2TCSGxM8NjBZC0NdVEmkzMycdL0BtBn64zRMuUaNYNstfNFef6qaw/UgpYhrs5
/wgm/q+bko84WdRU9bauev2J8RJxTvdFk5NFLtLFHbRXkRWMpv1RvdlbBmireYXwcEJFjJ0v4wrf
MGqTR+WPrlBeCH94GyBXZhU7SrR9Vvbc+G1MRnBa7ig+3puBX4LsqTmTQ9HYsAJaxmRvTaVTfcMz
EZnsOluUOugyVkhKatzvryVeawRCelxigIw/QtypkgxXq3Gc72zFCFpKdUNhRI/DAQIlW/4O9oqF
TSFRJvp4p0dndOhhUnrj59A9LKsk6BJgrFCbQfIDwqyeQje6NPCFkGs9nPjBsVkWU1X/XH9GY348
Ntlqcses/rMd+wQGBUBXnkt8C6cP4S3PWj4+z/7Jc40RC9fDrbfdaxqnboO8tmNUJdIoaH8mRJye
DZ5cSzTMbCA3xzmd8XCJrgrm72vX6lxJS470q9vxXkX2/U3QkVaYBiVZz0j9goGr6VkRo5SsXkTd
mbg0cfKy26vrft13nEID2/DrHIOzJUamSMEYpCvmbjaWKtuv35j8eMhru5cgFQBvieM9MYZPHJfk
zI3gVE4YZWjXUJfjNOk9EvnT5dyQxL0+PuPer5lENCFjijKTwpGml+Cfiv8mp3ty0UtnKtp1pEPl
NN07t/QGx77XBqzR91AJHWuQbRcju4D6Vx6af1xRqkoUVWs/OanUzK4BfwamT7E5MuRFII9MDsFR
H4hfExHuFjMVNz6pz2O4ohYpXSFpJHP3PFhwqn1L6xHRZwaDthHU5zQ9XNhjLmoN4a/4Z86OwCZA
nADcBj00GlUpacdJhoIby7eG5mMrDJ8aHgIV84Fh3nP/2NT6I8ws1tNK9x1mitF2CY0CEdClzCIk
6lUtiJ42uGoi1u495lk+yyyaTFa8a5+DtxtT4z/hLJgMzpPkzvwl7PBSzFH51NX2n8r9/SA18gOi
rQukccQTzt8Vu4zq+9SCKfwJNNwp2MsA67i+hHytohU6pIwgUF3bSI1fCkVWb7MhxPK23T8ZGrUv
tlfdBgAtK9icLsVxUq62Q5EYek7+hheH6k9/x7OOAPDS/bOlH143/PJFIcivPEteIVwQ+qkTp3yq
VOvyMWRAgxlAKXCeXQcv04aAumLmx8oOvPqbMBwAVy5xZNLYiIRfh3vOaVHJvA0HPyEmXwlmMfC0
Ivyx5Wd0iSVfjA3hdYC79fpbwYBM2VRb6LLEs6EFPGT5HUjlPuIoyLDMMdSSYc88W34hXEMyQ15c
/8W+lh9aYCMBvxOgA/7tNCqjtl1baibCJIJKFsQIK4NZwqv23BC9XghJHJ+PxGr2iRu9S/LEay7g
6hdbMCDkZNiCOQeAk9Ju5cowLmK8EbC7BvMiTt7kB/tv6kdnE+KH8rM+y0Ge19ZwvdssrFTTbiBh
LITZ4GiRp8tz0YhzSNNNd8sezCfQlQcuRcgVZ6TxzY2Wr5m1TtI3H2UyanPNeF6ziqqUcrOycVjF
tMuKBpcQayKtRGR2qWLYmGSu894HhVJGaWVhnEUBg954zINhaZcRmutq534F+XXO0Gk1rc9FhuFF
RsikDjLl/seNNOIiVcdSqbJaB3TEY8G9pYohR2VwX4FgpRnkKop38EerdtDfAfGtc91L0X+JjHGz
giyIIThqsMDZ4mi9NgN4R2PtxUENZMj1zgZqffTIB1BfLXRErIqjk1lgrx6kSptYUIER9MB05yue
PL3ObJkjSrT+IFrjzvPamZhHCaPCOl2+LYDqfxaiOR9Vt+1vQ+ZcvUBnZ4Z3yTnxOqhx9pSkxobl
siFRjiHgbiu8sTNgWlveL+rJjlnb0lc255f729zqOTt7nGOgrJvQoysibfBuN+cW2mVEXd0Q8KDj
2F//RiGfkrjKS4Zfja8IjAswJFBCvxpWwv5BkF+rocr21Ueunxi3I0n9gulxUD6YhLfYbwsppPGE
brKUQaeqXsaSJMuJ4bQAZqjd3f7vdd/vouwmFBUVUxZDT48b6d9n9eRgrT3gxJVU67x1KjQsYweA
4nXuw08aPKqNa2mJK9G+sfGaE/ZyXamHd3MLn0z+NCsKURbxOfsdCaUS0dlIEiO3BNDk+AEbnRdz
nIb+D83TZyorkbEH70ukbmZs8w7SyMR7DsBmzh9ppb4Ic8sVXzxXlcLFGhyx0nrVGHoYo+wa1WQ9
CQ75/EWYqFaQXWgqArgpM8dip5emZPV9Daq0O7SSQEQCDD55Gf9l//D9dB5cr//LmYUIgCpT/5qI
FFl4IEI196ELRRSqCsa/Y3TzSiAedTmTPqqK0jucedQf9MFwoH6NtQxeEheTZ8Yu0EG4nIg5Sf8c
IP2EC2JeF/UvCwXg18To2xe8sI08GuSq2SoQny6vNt1Aie0KZ1bA57vG/Av0K8Jc8ewXzr9pq9i0
istYyFYoT2XHw6g27vtubohOySwXO0hG3b7JxWCj0nqezorJ+Xgq5Xa+7kQ2B7JxnbE2AKkp6zIU
1xpMxCINf3Cpl1fkz3jgZlh2uKiZL/swiDvPokm3YwnKyQWJk2NvMEy/1VFIBb3XoOxuP9op/64O
OjLSaOReabgTkRP8u23tNqemPa1XxN9Zf8aIssxqL/FQayHTj+Lhj2/cbn5zcJ9+St0rXwDOFJdO
motO1fbJMG63OBnsohqCTOFuJXbb45k/rIhZgosmB1dECS6ME8TFYayqrxtfwFYMgYLOC9zMDW3i
f2xEM9+mNrUBM5TCb1pNJhHwndzVs3+s1YbSSgnKLrD+GgwTqMTuDlKrgpqi4/bGdyBAJ14yFPai
eTB1lVD+mf5rcaoPMXBMwvTZI1Vl0LL84Mze1mK3pVFXe4M1A0lJ3Lx2hyWGj5SKVR21hwMj2BiK
hKzXRDfa7Gz484T719F3uVGxOPrB29fsq3xDbAkqzkZMadEj38vY9M5lvMPOU0AiASkaQ7ebMhOV
9erkVj873n9q4kMd4UqT63GY/bX5qYL+or4eZbN24KFbe3RcUBDgvdvmlCe8bdw5hF7nd0u/1LcO
TREcEvUiEBuB45DAyuJumZ4s9GvebAojS1uBT+zRFTRV20hRs+I7UkEqq8/P9KMfKrltrZV2SDNf
dA3nHMhcXKYOiRC59uGLpVUnnSZoHkYKSFm2pY2slfg46Ifbwq6EdYBLFSftBWR1hiJhOo4laiwj
YKdw42CKZUt09hXvpObQgtxqmvhimPViGt8cysFfuUcESHwyuwJtCw2gm2Jq+mnX6LFffTXLJqhx
VoL4rEGuBAClrrGgyGUNJ6PSgRvrBBBy1tAl/HbuZLlTulg3HLKUKH5WrXpZkF5kkOCTkf2LXQ48
4+kVWcczOssQLLk3ld6xCqwx/TFGnLgRJL+xE3vjON7z6QOjI8PBzc7tp9tPevctOoEn/swQdwBO
lpfl9vC2W7ew6oaqltnRxK17YYmdei0xjWy7wf/zTXmjMTQSsy8oZ1GhDBTayDiiW3lHd0D1kjYw
kwH5aH/7vbYJsZ0qxZ0jU6nIax/tOO8UvX6I03KtmXdP90bxGeNzLhGPzv3f9txUTXj9+S2z6bEl
pOJRDgYhkGwvu5NQDqgV7Gk0U25MDMlz8LgYjijQulxE0jb4h1r3HaWBF0wWcaPoTZ4hXSGJBd+f
n4pjjQ0nS9JNMlqESasw0fwzU5D0KGckwIv1ZpVP2BZhEBxVmFHXSzbnhnuMHTqW72rzoghylYU/
MFaFJAvd/zU+KRTrjPcvCtigg0a9vMWj+IcK2xT4QBLVzJmV3Fky0BdqenCMJTg1BsJ8Q/sAiWy9
vXfCXBbkgqUr1jISaRO076GUwWcYPcX2/Kp8HlyXSFO+P+Fuy6bOLdC34NkjVNlbIYRICpBXBjA1
rtUB+2mB8mCOmwumiofQOM6X3PrnHFzzRiXVZGwUFrUpzWGND4ZkO6AGKw9JSfv9MyhATl2bG7b4
GX1T1yC1CYhMhUsxd5rO6Z3rD+1ny6ZYbK4s3bXi8OUP8L+z7DqxHnMqyPUb6mcdIF6yXZFSu/MR
w3/0BEr/hy2OnBnFaoVs0RA6ckM2mCuKrE2lLxVVQO1xPofDYw/YJi58H8KNn9flpMqeqEB+nHeZ
41ejlEIi+6IDUoWg6xhFLx7SuV13INoZ9eKUIkZKT0isyzbXJXRedj+TNRgZe2O6A1bZEBqInQi/
VOC7vbUnvwiYMGnq8USzn+if0Vnuy8aAVRk098vRuwr1RkH75P3o8v3+QpZGy/MvOE8fdKOQ81P1
LFJ/ZJ5XAeLQmvxAKK1mvwG1wn6LmHN+UWTDY6MRoV2aCIQvM9ASJBrqVZ+U5IYQW+Q5v0CcqcIw
paV/xyb4P5fIBZn2PXyaXyc9HtYb/KMT3ymgY0SgV36eaEf+NDmJxFIev04k9nSzPewHv8FHmSGR
+lRsbXA/RQR0j//cng1bHQALXM3iMtwjDEWyELggm66/UBTPw6ahM/CDqKbreKJSN0Zs6AyBg7ov
f0WM7JLd8aF07S/9vHeghngz3dLbDLH0rBhUg/7/HxkaNRzIbqRN1+y7NsXDzSUxxMNlF0T9XIGj
tV7K3/MYMBO/l3Fo6hZlGi4tr2byDkv2Q4oZLewSbL/Fp9xALbFlT2K42VL5ckLHLue0Yd2OfxT8
blC3lgUhzRh6dZs39pElSlPlS3G3RQKNXZ3WKCiOOe8Z/hKaALs+d8iNOOLfdEmxjw9QXfoKrNGX
ZvwuDkakSKDmQEwhklH7TeeWHnHH2J8AlI6FxI+Ltpd7gfjhhFtdRFSbUFLaRCVQJwhZegEdgPWu
mOfQN8L64Z2L1b3VIUScu50mHvjD/M0fLBJGNRvQDGBZYVdTYfAGDENGFTd3ieCD6l1ICqXou5EN
FRKLNWHvOGCIZ1Bc00R0Y/hvqoEkcfu70J07H4g+cYlnFrwpFVxzVp13HYJh5PitXy7iOf1yeQhJ
jYlAzcQw6zJDYZRmansbAeFvKowLTlJIokP/Kl4ouA9azEc30/dDLUtwUZ48NktREnXyt/Wv5uiH
gDOl0AzrzYNIYCmz2nsD4KwIGdorP6Ea+IGtUzJohpBmBkjLqe3XPtaP0J7aInthjqy56YLGYDNI
Dj09AtDWf6Uamw99o0NCUFxwgwX5HXMAvrN5rE90yzInZFeskm+4Ky9xccxQTVtmWFx6u0WgQPij
PbfodHPZUwGmV8QXtgVd6TeP78j17ylRVJ6M++X0sZWdXuiim6zsz9sHOXBf99rwldF1zjZ5yd7M
3VC0cYSd0nGriC6hQbCiEiDq3Jl6PFVmS+M6GveVBsekRN4GdkmGOWb/6MWlWEHOrdKFNGWcpKIc
pJt5zcPSl7fRWGTxaK7LuX7nLQX/XK/MvbkGgxXf/Q/Gxfrt7IRLOUfIuyP/C/ipXs2e80dr/7Ue
//9FlRq/OuFJMEij2jUUhIDm0t6cW27wGm7kNtlrIJu66UpJHN5cZwLSAmGA9NXFOahslg5a1y8K
JaisOSzvJAM4W/VTLxZteImyOy2pycTY30yaewsjYd1H5cziSKBfhnZtslo39k/ocMOLMAJcVuPG
nnXwBcUPqmVvNIiNGwXg6OBtyL1TzSm5MleK58vMwzehhO9usJwg/djtku0WYwFc+nZkkJpmJfUc
UHjZ15SpqL6aXG3YrhG3Cn3C9Rne3S+RxqlJ+kXVGJY5MMKMUl94FPhqrCaZti4rAm85WJ/lsKOc
qTIm8y6QTgWvdP8Zp8nbhTUvMgUpkq53Ele+eNelNbu7B+ojXMxFNBqyUZ33osK5NFAAzxETSv1a
36wUhkkTxL1Tmkq2SaY2WUMEL2XXSz0DXxTagKioJ2TV/0yvn2TNAWw4WynNLYkMksEId8Db0w+0
/YkejgqZztAn/Ygf9OwFSSD0DOOF8aSpesKIIVjdWZdReI8GgiEg5vk6CQ0+UEFkBGm0XAfdfzk7
vq99qGFuEpgf7kimikLRUwtFsgtHwfQTRHxml4Dr1/+C65s6T5wMMlGIQ9pN2+p2HOCF/nvVlPpU
loRSfAtvGmflUQT1YfGpPqdZzx9KSpg5ssP7q/A3Em/NP4b1GXQ9oFWNtTD4LczGqRSMpb30NZBz
QyFCD9eSuYLK9nanTVe0UbvbXIuq9bZLfXONSiGTIE9KcUe4dlO8yo8tslSw7Zbq2MW3lMGPZTHg
0vBiCCD0sGM3b4W6IFJHAmmXI35sn3w8zTfRD7OaeBF4J5FWHFTjRAOwk7NVeKOaSEegPSBEnSaB
Wzd++NEBzLVtsANyHAf3QJL3phUl7upk9FYESCg1yxZsAgpjc9CmF1kh7xwNVpwYrzIzqSGjPHwu
O4iMa31QDS1OPIE5mlgdBynbzfBd0yhQ2anyrK4VdG1ks37kYGw4HcwXv8hR3ufbXn17jdFhPHUF
6RoHkV3MsudLpDfzqlalqprFwEa0x9zNPMGVNSMuAzzygvifkwVj4lVTJIKWlkU6X98bSi7Xbw3g
KL7F4BuRA6/FZDS8UK1wY/CdmccOi1NJ6kyQMPr7YB8QXHuBzGKrqUgOmCyYPrC5Dy4NUPqawazb
GIKzkcI6vH+h5qv8H7r8uXXNqKY72SssSqHiQwaw/X8RgoMHbG4ES4QUG5gZqJWge8nQz1obPX8d
jkeXkiC50gmtaZbSQfJP40x+rYDFZvjkKtQB2rBXMtCklTpJ8q3bv55JTCVQKx7OcZUDlUdqhvB5
R9REPEHKjRodQoKl4Rh27Gq10cqgDQMRyGizLMfQPjKQTMSsJrr0rHnNnG37RavxAXXW1WI24Pk1
nLFJnumxG24I5O4H4o0A4rVWgxxUGewLpYt/IEI6EiRhbulwsIw5rGdhdVWELh/x7xC4GLJco0St
nVW03iuEpZiuPVe6bx9Inv6iXwvylDZHF3x0jyWOYVJLa5zJJT1sTgaa9KgsnRyR44gTiyw5YTbq
/QqsrRQ+NAYKYlRHt5QzrP3jh7FoJ+alyYYSpZMu9Lyra4ccRX1rWSK84owA3+UylFnKgJwjF5SX
gBNF2Mgmh8R/c4ycr6oL8Am8ikirDcKtuwk4VmJfROOHWEbQEEkn10vjDZIpDUk6ANtA8w7ZedM7
+8l5LIdcWE46J6dGXQ4sL1MlEgNlwjBe80tq6G7YvjGTv6/0tzm0xBBrzEvqIDuv57NQwUjebYHx
yxzMOPiSdWW4evRyRdn2AOtE+1gbIgbNY+Do/V64TAolBTvi+8BswctxG7tvZa2vRw1vwIEgwF3b
JPtryjh8zBYnaOyffm1ggOlf3GGVHr8FfV00bF1gZZoxyy8IooQFsedt3dR2PMTk6hd2UE/s5IDg
b5WFMc9dJIfB3q0cMKB7qnyMwF/IfVi42tPAhnwX699awIo+dGErgqnofSFp4u0gJ+GhznNDtQVL
GHmtwBpYZkZu6J3foY9OrIkPW4ZCSwoLL1jx969QHu7BYJtUnOSB9Nw85e6LG9Hmc/lv6LJKV+Vf
V7Vo3QF5m4QQTTuoHM7pNDVD15g1Uxr5uSyE8WnVF5KnKOoOFKh6/gSQcKmTg74H1FFiKv+skiIa
hNrpEYI00tTMTXLdy9xKcva3jUxkhFFj2FUX11ltn2OhcXLCbLBSBY4i35pzsw1h52NEiQMEg5ya
pydjNHuKI4BG8BRjLLfKc3/AgG94rvHeEnQmIN7cJzer29Ojlfs0KyPkfT991IM5cdc8GNcNnkxx
K0gOteU0i09J2Ap6jqqfF3sbz7914UyWfoP9xGMMBUFjwe4Y7oayKzhX6DGT7CKpLyHyTd3k5LFZ
4m2lNiChEXIZJxNjP1+SP4z10Dx9LrL8i80vOdvCu9foiw3cmCtick+u3iaw1GBdRiFHOfNCaBX4
EAQ7aWQ8Dl74Qy/5jeMA9mlLcTaulcH0uMDOKF5fWrsFp4YCddXgnlJ7mi5lGwZ+g05zJU0cnjnu
vtIY6rC7O2Q7hslsud4GgWQU9GJCoYfZtOcqIObv98NwPWNgwWGK96P8xz6oVYOwApG2uOcHfyLb
NDbI0rDx6R2rM0asO1jFQ8JaOc+1oAT7Ffc5CjcEOw/PvW/uUfqS33jEpJ8yC2pb71fMzjxYR0ui
oqceN3QAF7sBNe0tFhUk2zHlBi+CGQdSPrXi27Gl8vz8nj6j9faOw0NRT+yOmxh/LwxnLN3XYOFp
LmTQSTR2zV7COyXcDz6k02TGu+ilWCKNyVBryD3hzxc1jgzj5YePBqwPm0lYmB3DTElLVn2pCt3L
rSmGBUIBqzwW5jC46Mbeplvg7T+kV9fEJLSWf4AMbcY8cQYLRuDWXdUhwVoG0s6TKcEuHRex5BNG
6+7YJeXkcNhoDq8Vyf54yAsliNj162XXW6FliIcg9bOLTAHszVUreqCDsqizerXa2NbBWVGBeI4+
X6vGoZSK4soCOKry31UhqbGGd9uUZesQLk85XczKrKhJbDq3AfPzPQG64gTCgqtcAStvdHcWPOAg
DQk1Wca0iiDgtYDPFTgAGk+9zDkKq5wgWEY+b6q7quysAvcQAhg0vIpTTmgYjFfMjKfFFMxcHzkC
76AUNR/WC0o6cYUyqrwp0eUFqQ1w15Re9rDcv8ZlWQUyqkIyzjrIemTkSJ6ASQf8D7/SusmcBLBn
gxqi8s70uCAbRxv5xRtFcojpKo8e1RPMke2v/Hp+2DN84ECjCx0CnDuMi2b+rUZvVlbapbqvGsUx
BWJodczzvmPcSMBpqaw+a5fL5pkZ/atWpAoXk92bFiXWLmgjq8nCsxci1UU45YZKTYi+rw5W/8/8
nZcBBn+pBp/t10PqMQmYGjdbfvMrZ0gu+Bd91IUt0HINadCpH93ckZu6BaOPoVV2N95AVHEoGJiU
i6vJLAdJAW53zb9kdCfbIJZ+JUJOUXCPuvHd8ciZsUe+jPh5H1mWUXrpaCiewhTjN9+65ti/Er0c
DqXUgPTOk/eUldvqQmM+nipTdJBe/GO1NDjj86I8ZeJsuJhuQ9x8GkqWptqnn4l7ngLyJF70BX27
tgfWNmo49NLti7wR+BFUGlJTObkvRP5+ANr5z6RKP+he0fhoomhgeNQsly08hK3i9HGoCC2hp7eo
f6K+39GOxnB/6ME9CITMFa6wEpojjQZheUGpIp65KmJ4+cIA44CUTQTXoAkCgEE7ZknU1OFrol5G
1Q3jgnw2f86ds48GKGPinCn0oRWX24L20KfObVi/q9cyx/Mljv4Y2yfkUppMalCJCXBfPt7nUnQY
cZJCNlY20hD+1gt5PNjLy3QXfboQ2pLMlAJRnUn3cvMRddLFL9bw09rF1qAopd80rb9/Y0zWLTw6
eMidoJz/GC+HUxpC2WnD5KryX40fOOaQqnn+bovbDjrVbfEy1nvYkB/tYC7pZ6bfAVfL7R+PV2Rq
u21pGGvYIMvS4xEOvurG//jbj0SFvIzdjyublXsxHI0lReRD/fiIseGQahJlzunCXgAfUqgiCPua
kjswIy+wdkniZ53/ESr64TZJuTt4AH0XFKDYAQyGKAb8mUD4/CGg70Ntsgau+7TJyeteyiVkOioo
b16a47ggqPhKtR8+uNdo/W/CHmGNmig96biPFJQUX4NmDAhm7t+sYIR4hCmtGePAFg1Es1dfc1Q6
DFlXKi3QYT5O3vM/bHPQJyhZ39EopW5k73NJaM/Sqeeuq+wwY3arFbBMywZnvWIwNJ523jBtDWnk
e5kOM8vnl09AcDESpPa60+kk8AtwvnCrAl8y4vLpX42A/pgGguEzPr5qJZYSuKHA86x3S3VdjhN4
ZHElbYaJKxfZeoMYZQzsNTQHAVHDGG/AGcLfgyy0gszYxb6FDBR2Hx2ewyLMnBELhZDze50rz1uM
Z3R7lux8bQb5lOV6JqZH9A4TeWY5pIxV0hJOO5b6SQhD6xc6wMl4Y91z7G2I5SKx+UxwXjAigzdm
eiwo/i5lAAO6o95u5JoCeZ1WhmvnJu/p3D9aLryZ6JuwyUM4SNSlbn1B6y7HFWXNv7418covkELt
gJDNWtNAK2YMdOl8BxkMe8sazRUeX41hEztF9waRtu/4DGGm811P625lRoR55fcEASfbAW0j1hPH
LOeAdeQT0Kz/e68LrILHVt6atFsCiklZ1M6I6L05J9OOco+kaxJeeHQrIQWsRGEKixvuUjPMEYWJ
AV3qCtZU3a+m7N9DXBGCpceRIHxRqArgbyEfZq/zidmJEdrx75TSOYIpuXuld/XoVHY+emGB+BZY
HH3FNwGWWuoppq4N++qeMqvJHRyDVesUk4i64d3iiVAonBdqSo8W48Fu+aIW4lZFs+wsaHIkuVb5
DAvBPzJK16kMsU+mkwAS2o3pKsUpAwgdsEcGZPkmYjACC+Svd2lF23uJnD0dDGm0M9shVmJvJUCj
B9HknzvQU15SNbALGNBIPj6XJyuhSFcgRj/c+KFG6lqoWxYpNjCq3LnVGuU2rUsQBHKsjapj63Jq
d4+IH7+u0HiXUFVWlheIbppRHyHqd0no0EqHJRj/40QW/c68o1Zogx9MJLwrUx/mQwhVkyUhz3Oc
AEsCAUd1aZon+Xm8U2stz5T3hoanZ/l0dwNflu0gG4LmtS1HHxBVeHceepgBtns05NTT82YkylNn
NeK8yqFA76+82p8DkQDVRM7iMDiS7zdMRa6Lf+n99O2sJuaQBN2m9QXdBQva8fHLdnx0Q5+hEda7
XOV2O5gJVr0EhrAm0CHOOUXrDqr4GvvPqLNsIgOTo0hfRWwed1xZn0X7mahCGrLGcMDsape7VXY8
ygSm+pbjcES5vfDUNHevEetnJmrJwmnmG7BIRgERbk1zhLXCFI9KCyalhNHrBiFKv4X08XMfZEYH
kignsYcAeegSJVA4w/RGkbBUh3vShFXQDINUygPv8/0+1p2hwfxFx+iUbgkuWMkxZEYHNsxp7OWO
ND0k7LdI031iTSpp7/OeA/fw+IaIkAuch9Gya6gqcZKy7ZgXmyLEiTzbCkt4xwwMicXoiJ/DNaCV
tgDLWgKFENWU4Zikf1RiQLmdjg6/6jSWOrpWUIBk2ZVOw3mgWOYsMQVtUWYHGYdGVFEKvesaqsxl
OSeYtv9bcVDtalb43k3WpVNgiBWe5D1gtJdSU3TfVWdm1pSypMywzxH2lvLtL0i0dlBp0BVQezUe
k9xiUF7798D410/VVyeToDEC4e0FoHM3n52JQSIfnPbjpzZP155OQoUn0vqOx7KU+bUZu30yhsLb
nAC+ssR1FuqpYB5dpfw/qHc+6okyRV09wuWF0Jk6Ea/DspN8hzdU3vZjUPNhcR4VuAWjKMWtrJ8K
stlzpw48AMhQyG8FQPD+tFnxzruHtocOu2yrygscuGk1ASa605Idf8JlN32r5yT16z8wMvLWuFOl
9jw9DB4fUBYpOUmDG9J+3hs/h0l4+HXOeLtOuV5Wncl8mnklHlLH8NiJxZQ30iRlWbNbvSqVNkLB
xyFG3lRdsyeYfa0yYGRBbckQus7+aQGjG67iCSWUqZGPXAzfjHbN5ZwNiBlIc/KL7nP8i4brYL/0
VNxsF29/1Zhu7SE4yl1UdVOixoRjKgi1BRYebrwFHnJSla2Oqi4VnCmRzXVg7+RmmXody/hcbi18
OS/QWqSOM9rB8N3brjkm+6+OkgyTXhEpiTnO9MCsBLYifvweQ9hYcus+hpJkSzBuev230dNybBIR
DlFhJuJZHMlO2AAjr+nCgHvfAJvv+KpW06iLjfY67U88I3VFk7+blVDOjDyN7kKLAoYomDLvNhp/
TGjhGWubsHNUnyi82JQxxer0g+qHpiIVzPA7sB1nlHrJQk2hTlGSwNYE2NkTAv6yevemUDyWZJZF
0H6GOqe5dLEB7DnCNEI5sQBv/GDWsc82+WCsplsgOiE9YEs3NnD5VaVPJpblyZEiWemIkwOO+Wwm
otGVML3yrg9tEkRWSSoSOxRMl6jdR3Xha1wGa1Rkc5+hq84AI29Y+19DN5ATUSTay4ZvUUaYHF5N
nh6BIEF9r//CYsqNhAdGCifrrWxGAuUNC5K+t0yfxPzYevMN0CSLvu8EH5lQsJ79K9DHMarz/DI5
u/t1MGywLldZER8kOkcMdcU6p1M6INFdfYWtogy1/xBkA5Bykhxg4W2lpQmfvtiiNSZWmAv1ttNI
wWpvFImZKQGJhzgmTXCFD1DZukXRre9/T50ullEf2OwClVLf0K05goZO+nwLiW69N+GppkJXHlXL
BmDHe0bPZi7WssBUc+LDEpSw6O3OZvak9b2RIlosxPsIEP+tP/IoiX2BBjk8DvUTTgTVTSZ1oyKf
S3JKifi4gX8WalFFs2Ugo00jlSWvb21ee0MkJ6+MnLf7+OMmIi24uBoZs4ec8pGtj0zLvBRBHv8D
s9PMPAybEbrzynbGXwkQkBVstTswQQWUVWLSESxveWvs2SAIGsCv6crpzwRgsmYupYpVHlFRrO8W
fc3qcBj/BrcTp4S8BN1mMM4gzUkl1og277ItVfUu4S3/EildDLVzPoqDx5A+vU3C8XJZnkxPKAL1
Ys13rtpXMu+MTOT8zcqlR2xk1llPvlf2lhsQYi0KFLVlBkRAWqmhdbUeuUhGFnX+hSXDchWH+vbU
TThyRA0pF2ly+NLSyQ5W/Mf3JlmSYmoaWn0qcjdTWKubf/OY4N1CnNpDUjjsXFFq/qIc5h3zsYG/
Lg5AbbmtKd4EpqVX/8CRz4zvnbBWLxCcO0HYiuDbZkSIujirK3FL3i71QzY+l5Sf12RtksMQEkM9
sgw56v8qy1yG0ma/A0QsFKptAdTi1kDuY4RFSy7fg2W1qtih1A4jU2tySD/2KF17wgVSDMvBnxv/
f3EPGUz4K+I3yBWPpDCUZFrMI6SmHJd56ZXoOkrgq2LaOEstz1QmcwtjG04C0L8ok9cg1pgrfagt
PH33vViCiZDqGfvWRNdNRAhRyFz1bIkomjGLGTFgrxs2gFZWti4PTYA2NogoRgtXM5BAzgxYq4oT
cLOIDcxrU4KnkVjCH/b1DWhi7/+6IYTFHgpKIbiXWXcoApsyNY6i4DYqhokv7ZUTW7GEvZfiD6+x
lcS5sf2qvePOkapNSIwydYSHaBOYePgl7USmGX4gSP8raQoBYUSmXk44GEVmaEETYug+4EcLTbT2
5MUJno0Bq7r/kE+bHw/iNQuJRC02V0Jd/MBlIRMCNqDnu1IDksGIBMHCn7YKyRVCop9Zjy016V1/
fsZOZr+zP9ik0DrXSynpLUy7sMosvLPv1IOQgBXdW1Wallapl17eotn1wQkqKm5Vk0p7qBRwsR+i
wUxOhc7IzcVm8B8wCpDvVImvnCFYNWiHyEsTjxwdA1mEBHv+0VzPI9GjJpaI5e1AabjIXKq4nM5z
dpk5U11O6ryjU+pJLxd2MvRLp8i1J0W+aabWwFj8eZEo2QLlIlv4R9YG4/AvO/Pfj/tL3Kfp4yxn
xUXZBoOzOeb86xQ3Moru9WTr9SGImmQSk8ZiwL69HrmDT6YBgl9etFzhYZz/qigpO2USwHCR0yPZ
u92Z1hwdvMUfyiNkr04980yEFN3ONum3r9tbuwGa/JRRaJfUeSE7c70F3UN9bGGsk4vKx6YohQ1n
yR7uJX7/jaYYAcjzaP2YyGmLEuPaLwI/dMee3dKDA0mNJ0XUO4a2DKr3bGhaAF71gUJNWJ5/Plxv
CeD/Lf3IsfLgX94EQvQhoA6HA3NPtp4ZJStZr2L+DIs3/nNHkoW8OIkt1BWxVZPmdiTpV5xTdZj/
uB6Ih7AqApy2/KvMB0JyX7wmq83jVMo6frZVKLmEeM0m2Z2DwYKMxOF70ZCeRjQL8cXS7rSo63fX
Lr0PhuKh/1PEEJUGEdOaGg89OODh+yffXwR72RcYfZws99v/pI5SUi5Ez190Y+NqXoW7Lp6+fXRc
f8/Kz/KvoXY3teSMkT5D2c4o+n6on2DMFVDRoKcdM5gLsugTwd7A5BzsGeHrwyDKDYhFYPhytFTL
9lrPsSzhZlk7Gr0fsXEgYDJfO4GggoiphvbZHfFbG2vgszZqA5uGySfew0SYOx0ArVtJ4VbX+HHV
EQXMk9Ugss50GzNf7QFaOukKAyBQbK0lFN+XDAH5aGnu1mNi0RrbYliva9WQyaN4T6o3YzcNO1DU
UF0+a5ceDOncmJlDaSOSd+aIc/GMpWIphodYuUonKC3C0Eig6lhFBN1EulIBfW4z2lW0vHZP/NMN
1YzTz6ymgbl4ulEDJ3C4cJkjjGLdl7nJCP+uiW8UD5Kk3wL5lTrrKYRiuohER3c49FcZ3VFRKkul
29G/gCPe8FPAfjLxoMtbuafV9CBBViXsvOtkIBDBjHMpt9veEKNZgj7t6e+bXB6oQlxARnu0Y8UK
T9O/NaYJeXJ9oXhnEAFVumnr03oUzO8Ym6G3YJFF+jSRLogOxiK/5juUAKE8T8xi4Jxfeia2FU7p
t8zyxxCyl+9zh9pxDsBrICnLsgSbEMw1MKDSYzZl+3JfjwME27qDGLFeTydVh+kypAgbGT3PefMZ
oPNqkzGB93ZWjIQjBFY+BMUB+pxv01zQf/wqotqWupZ6x/k/r3yRXyYBNCRSjwqNMPqDT+/eUflQ
+ducdXXNHIwXwDwM2/Bb6NXiW8NBxS1V2lWlQ8dpUadY+yGXDTCCwlxmhZAzj1zrykS6lJYZvxM4
muooMoNMt6IIEeq1Wl5zC3i8NRKt5KS1dgsSOvBlWR58ESWfaTLqcnasy1P03GFxe/QVm85ojcCo
FQT+++jMAuITEdsu1pDlzbHjbugCAS+NYKIbnUyd+VpCqIydmTawLeBXPgZWui0wv0z28qKYA7ss
SlZpR8wlPdO9NUn3nrGVkfhM5mQHN8oM7OzGMlG1CsVT95Ip+6M/LwuCgWITBBzQZkQKX1bagfow
VwDUM5kFKV49Gt+6he4Q6OQ6dyeAxmJuGasONTVP74ELFQXgSw1DKTE3ke3PdWsrwS/ZnCeB4LIJ
Su0Wl1nfgCr7+zykaCCNf9kesMjvBTe+isGFzM7ZkNn2So1mK6V4XoeEFwOBgwZiZPUiS9iBmoIU
SJQMyIxiYiOhMRyDgARFwHYruxP/Qy6n4wSk5mKcRBckXwwi9funt+OuatNCfizrkyKwpysRIoeC
ndKd0Z7yhzzSgrqUcJG5qu/xS/6sOORgwUcjn4Bc8fg4k5qccyC/5xCbh/eVaTkUFETf3K8R13Cp
0dKZE6Rl0DjgeeJHQCfrG5LFyPTIiKGO2pywQ9lKNK2CrE6FAU2F+RsIKp35oMXrk+IJW26/LExm
WdggKq5KX4yBtgK5j55Re3D9SuIY9eCUB0kQ/BWThcAIac2GWqJj816RDaw2qaijFpMFi3JY2sbS
6sC8FsX8cg2Farya6lSQTDWvCPdeolg6Krk/7dnDG23fulBkyRRoQOuZSTgFMCWTwqde2IeW9HwV
U30kLR5vGir6jSVl2LPMOskyEGa20u8LiAggsOM3geljgVNyNYceUZgWgreK34lH0otoxYINSGxE
76DiwnR2bpQqSX7bSgZrJOa3UHF7P+m4yAhjKuuhwvqsU/9hXyfWFOiaV0dQcL7Sl9/DX8NNlbsi
+2GFLGfUmglsENAZZtLQYkZLxl34wJP9TmasO7ISTYw8CWpErdmk3x8hEA/C4NqmT0OILSSdnm0b
6BGtLsHNa/pMiv4ppnGYOX3l84Z+LtcmccFJ7mX4BK/2onASN+ps4g6t6OrGR6eksTUWF4ymMye9
vTgiLOP+FXcXpKXN+TOWxWDMXtTaVqbmK6NI3Q6vxkmyAY44Sc87uR6CP4o9wweelvWE/32dyT9w
p8AikuyhNxJrOdfSH3bh5uQYrpRT58cMjvFLJlsp5U1HkL9dplo5nfbjZX3ua3L8fm41OKldFzUZ
L3vuJ3USSlH2w7ZOVD8t3oyEkmeTwtg25aNgLJFq+p7y70p41HzMg3wMX+//y2g2JrzzG9I7ZGvJ
3K5bHy85oU5wKxxxCuiNvnXP/ueE/nlgpfsJi0E8bdfVa/p0yyWIiWSjOmXESxLwGFnJSqMxjN0w
d1oeD3V2IvtN+ndlf8kO6+8mJCqams5nJ7L0JarHhgc5dM8WLl50rrmSjb7Wo6dmI9w+hje3Wjle
DpwzULp4E+wazcgyJu+GhK8y0RbTZa3FghhETASJ/E+rGFLF5IWzedSGkXcas9kfzD9V9jYHdUzR
q9PzhhgEq8qkxqaSvNnz4XhU2ap1Ib4bJIYb1GE9mG+YA+1CYShh38hvwut4LMUdGjVhreEY/ua/
M5ln7ZskcNJZiMPb70r+gvAOPkKFqOHndcTy+abmezVEkdGGG4T6bkVEH4Vx8RRUJXhbdW6al0wg
J6JPOjgUAHeS/GIq58/p2b5HnaRR4IJCNMPGqssshkLXUKorREZgTZwa4Jwaov9KhgtLUf7cncb7
qKIKEVM8HI+93Q8i5UGQb1rkAJCir+jzpO2iIEeg/2vHhxEwQ4x3zJB4Ysgpc71tsJxwT3c1O7XE
zCYgVctGTjrxTvKlTKIkPovu6fquFfdNckUVvDL8QPCafL8ks2Oci6Pg2keidtxhcJtnnibWaPKQ
kCg1DHnBB+0vNZdbAto6J62nan4Zhs/sK9rMvh4rqeaDnzx2Wdv3bdkwUQugZpg74jtThFH9yHu5
fFXiozashrziPzDu9NjPc+0FZQ3rQzU8/l++nLUXPWtspb3+HC9Xq00QRrMEKOfK0/JpzWU4P5dM
Civ+Em+OlwNBuTuYwKvYjwqBwytx+Oz4+/c1aF+akUU+ohyVtLvqxVp/1MU2j5HeRT9nyHWYZUA2
oAIjEFQJgYDdigXmUimFueKtTaVEFn4Mhy2W4fWY4XszN+MBfA+PZEjcnwfU0tWZotj/Fcn6ym+o
N6EopSqn9px90bH1F2qtjLrL1uJTzEfadpy8i7REbUH6p7ePOcLam/acBLatwj7eRECYzgqXP75g
9CvkxZ9tNBefB1nX5dAu3L/SJkXOpIIjphfHLXD+wm6OgpEcgahfLg4NqrsGJGqtaTXs7kHHZE4S
BDUDwDa82ti+/Joli/mvCBmOzdR73+OZ+cLD2SVELtahwGRnii9kGjBXUaAnCQzivyBLIKCBbXPV
UjIkcrxHoPAsOmzkap5uNW09RaaMqRccSqs2M8LIlmn1nGdkR+VIinbhmfbKoqVoXRIXXTzpNTDU
8DrzRrfAE0ZjN/ejtQcVg4v100pphJilZ3avoaWe59HU5hUE5yEkCETI+jz4rPwwREeKa2oiegzP
6zB71prvDhwzL2B/SotC6VH9d4xnnbKgdVqRpjCBwk3Ug1ZHFbTP/WHpgqWKpHkp1xZZe3oPxluD
tstISWUJKys6Kf0qvfJJZta99dfV/IjoF9LsCTYOBHAx+IVHikC4PAVXZmAJG9Xk2DJfnNE1brnQ
jM3kgz/fmOwEv3EObmYBIM/i6Q3JcEUSHGmtj4XGCnAUv1YBVEOrsmbVQXbMmawyJ6MGLia0HGGM
E0e+Y6sDszX13cuS2SZU938d2sM9iy3E5q/BDfgWEm8UR3rKh7ovj8SDVCyhepO68UTwdSFAfARx
StzjHkmAgIg6gBO+9nkMNwdCd1j65wVxrBgBD5Ge+UIhXA2sAK/V2BMXLHZjK+QqvNN2oDhVrWlU
d0WiVJ/d+6yo1rCdeIOaPkVcsyPGP41Zoxj1YgWOaoZLskbO5xj8hI6NYTnQeCuk0g5GecCoLxp1
U6shrfFx/RDN2AX4fB8aZcCWOpCJn7QsT13sJn29Bl1go5YN1tKVdsM7uSp4g8PRPp1b2zEuX2OH
+mMzUFu3FWNUsR8CMUof/Oa2HBrb6uBELMSV44EJ2hcnG5CFDg6Rm21d1DubXLOSz6Q8SukxDfeI
yJ0Yz5s0FEZvDPEUBmMQ3QiGrpdClSJ4hnGSkwtBE7IaogBldBa3a9GlqcN3MHcyih4mVi2a0y6j
38JHx2p58j5bOFdaBcwCXa/F+fYNx4AgNXQkIUjD5ubudlUEWNR2I4W4+t7sC0Gl+aeUpy0LS0sP
R33lwE4lZ9jLOmwu32bSjS8ERCiCYtB0UPZ7j7DomDH2Jezg+vVQCL19wpir1ZvDewlh8oja29Xh
XiwlMSOznwSHbPCUx5B+nsoq/eTKWVlTSKs37UkSM8wIGzIoN7Gv2cwFbP1vwP/n7ZWW+KTubfsi
ddQwsxphZReeszvr3oc2hRDqQz5ESdjt5/0o/GsWuql0J4Z52CxhKrj2Q5b6Coc9XjmS4EfmdsVF
zd8o7B6Y74C2iJVcjsAazVw/dvUE08XtTfdKxkKbjfbqIyzU1YgUgI3XDJu8TTymfisEcc0LXY5V
yhTo56ktSlZ790efpjwwvBnccBP8wWWzGjqjFCdOsscYryAs3z/addDnRbIQNcm61UpnlzsaCp4D
G97IhUjnv+HQc4jKMwJzgsPjMkyXJkhxtH7SCIyHmuKir+Yl5NHKBCyAPCsO1Vfl02JwZ3UbSWq6
27WLTtXrLCuyAeRBcRpNceaWdf/36lC+95RyykFQVboEzB0GsdAJeGnkRRH0iLJrERS1iEzaBPC2
MTva1qxKKByki5EckkI+J2Lv85GQJ13ftdFlUbtfJFUJ9zNgruLz+OsEQsmGknn+ORxwFMyTL3vV
gld8Ba846fbgfURgUGjyLq98OUW0Pv1pL10eX+kWaiK0SziWmCkQGBJ4LTR5f0NW/uN3tkflIvjq
hKmRL6tYRT6Dv0usJNMM4L4FFycMl1FXiQ8aH8Nrq6NlLt/CIWp6wzx5+Aem2gnrdRsJOv7JG4s9
d+zXQm4AwgF5YaisG/tZM1GSz/4jvYQFLJXHYWbQ3pbZczGxFXZhiGUY+oyAHScHUDc65iv6icLJ
nSQMNvATECnXpGmR9k0Xhpcioh3TtORLZnNddCaiumWraNKqtwYrf8tjs+8EHuw9W3YW+6d+t83f
1jyXdSVEzMd/nMqw1XPghIwPATlnotnYyX5HLkR3QjcDmftQfStUw+tSIbEnsEIMXLFoaZzg8eUl
AV0Np2eD6W7GwIq8yANzvDwaDyi+hI1aaD8i4GX/KsXQyqAqKFviOxk+DXD4Cc+awkeMS0VF9LMM
0buoUxwehvVELqC+Cwio6Y5/YnPhJYHfh7veVdyMLItWQmW988IdQlMo0Tcc14mkxaoCLbOj7eBg
ZhbKgCovHHb5nGA9YdQsXYlx0+kFUU/N0ldJiw48urIGMl3H83cXzAcPuIzoetxv/hNOdE0caymn
Gbl9KCRRyk1VLRvc5J0ddg49nVAvgX9WpBAHm/GA1iw9pP7JZmcNrf0hSBUmSAqbWYcXrJWsBRJ5
VMrtbizgSXzY4PMCnfLYLhh2yb7uUeB5sST/ZeGzBKPRCDgJiB1eBi1/2/EPHgMsaVwKEEufLebA
hbHPQP0SzX9SgRRS7wRZP+sK67SGgdf4klUCQgZrLevORI6bA9WGwWqZx/bRB2iOMSPZRYRrYWxX
KgTSre5WUc49DC2XFm21+ZphjpRITqFQGD+zFd+rlyNXlgz038PZwwc7y9tL5ejtUeBFkJizrWgZ
n/3LxkicKzDx5vpyXnsoqu3E2JgEwvRp79fKh6Aks6lQJBZd8ncjoB71tnPUWrnuotVvh68Y3PaC
DsnKJv8wq01HJI3TRzBr0Kl8VVhOeBK0diXSmZb4CaHm1w00eNcl0l++RKK1RaU960TM8QWStqb8
VxhECE/+cle8rgGQjD23wjuHkFw9/MZsOoWu16vIcv7ViM+pfo3kw8d7Q3vGXjpkryjrvD8y83nQ
bqhDA8vo0+ZbROKAY7yfoSRmMOfKZNZsObN1pdooP6crSmX6PvR49vwR8jULZrr9Nzf6L5elwByS
SL5M9ka65zyz/HLA3xiieBLcpA9l0GLUPl1LOW34o13JKaZJyvZbOuLjbxfHkLF1QWH2nTYQoIUN
FlTATJT5nqxEnjD5tXACbY0Epf8ALtMxRtK2vEu67SlEzcS8xALv2+UJR+QYSKnYe0qrQdlQJsxw
5qtB5IJqeb+sUAkKVkDtw0dORpE5fkgFY9zaqsJtmLEtLqYp7pM5KxQFwUuPw5+0eYTjzz4aUxy0
3zYbLhP/QcwqkrxP/RORuuSHoa5h7H6rUgO+3ngDZQaApB8AO4zpJZ6Y22/B5KnpUMcK9Vwit6Aj
bmt5vW2/LF0mcgJ7RWggcaInsgDJde8VWBbJt7e3UE3ajk7uCHGt8ETm1BPETB0e0y1dJhlMEhHQ
u35KWcpA50NOwCqRhBe6+fnVTr/h6q1gc44EqsCzwBtcqJ1iD9lPMa22lMaV3yHOczX8b8LN6UJM
UX/t/6RtCn1UZgWIIfzNSlJleuqPtSsv5686aLcg1d5fSjdM108YIPcar8ZbSlQTSa6Ts1YSTMfe
sO68DvGM1G4cjAbmqDIV2qNPm+WsKJLU15lbzc9l/rb3Ws8VLWNu0/6GJv0aKOyS0DXQPDT7a9fc
iKpYA/pNy+rrrdsOzWgDmpSQVQMc5vB2p0tBsrmQxWtpoqf+G/ms+PvByg4AA2xZ8secT+huaDXs
L9f5wU0+JDLnt44jQiNhwzWct/kqPqZ81VO024bkPSYbRQ29MoK7NdFVktkrKB0mSsLVm3OnEYQ5
THJpIAkB4ozeY1ez4aPywGmkSzNWItQ7RZAjcRj8bPjbyJAqTPXqzLgNnNuDbq083e1/kZZOYgAs
trW4bveXOvQLKuizZGjlgfL10vFmTz74Ot0KF0Jt6WwFxOa5+ACCHQnE9vxeV8KOjSsFONp1qVmB
7BYtWKsK3AhwuOw4GcOhAAm3vV+ebESy95GGcG1pCVaH+M+C8IJu7bnja6+X9ADcu0c7DbMAczaF
pmEJ6v7qmjQeyDilGjIu3Jk/K4FTLd1jHP0yrVe8kHO3cvMq0dg7dZWFKDFZC/Af8V0rf4vPdlfC
qHkLpYnN+00ZyBbR8YH7FlZKN7ryR26wa+uDh3BLLq5Me7748jqvl7GaSMFpJ8mVxBSmPDASr6XC
I44hpmFD5zf/WAOOeeN4QJdZ6n3xX1tRRxDG4pAIOERmO1o1OuD2Zbh9nAmLahIw9eXFq/jZOF3M
OiC5OFgFxYLyfXiq9SLKg7cfnzBFQLk3zigNin0RQ4Wj+Rdtv2gQraS+YMJ7oNP0pmcrSpl8GAL6
ZB6B3H17GU6leP/i4C1R/WTeQEMAl2+KNjAzJihvAwJs8WvtC9sBn9vvouAhjQBuRxO7Nb/NDgtj
2NN+UkeKfppk6aJ0RF6HHJ94ZVp4CitaFPHp/Cr0Y6vrb3mTtc0ltJkw+DVf8OwBH7cHY/WPMDnb
s7SZgB44MDMDbFLf8SiRj0G8CF0BzekCiNUpPfFwQtpUWl3SHdkkInPVxPtfjQ4hrf2v+C7pvPcg
E5CiW8rexjlOku/yCOnrPSCjiicglSJOti9lWbWiH1A0fCRuQyTHWLfxIY64MEtcPz0/FkSTTkWX
LCn7wZFBopOSWFjM6LoTbdTHUygFN3/aAtEXII1pq22d2Q/4U4vRGMBGOzbGwrVWKh9l0fUbOQzd
vs8kb9FTm2fuMaVVtWQUQzfrNGj8d3Vw5fWbeqeVGQHGf4wUkWY0xnaKhs4n00fZ9axoOusDwSw3
xPAq7Iq1FrkLuiy9xvkbvGarKTX+gqFWE5pfaHjUla7h99Hgi9zSpeJNJzMymXYpJlCLTux8TNIn
kk2A0v9nvAl/cjmjtBHsa2b0DV+iewkxEO1VykvEPW5l8rnk7aTU+t0q2YpRDK5q4M4Q9b443fw0
5/xt7BqKkQV62DYNLVIpZQD3JHC0uVIipemh14Bb8jFn0vKIWS/AEwzHAzlMeO/H3mrkj58d6NmJ
6A5gq343AHBZzvYZzGjv/A5LW9x5QLYUNEB5nqD+hwnrMbt3UEiC4Qzw+W+qKSvB2CKUfjaVe5sA
4OGZoIzVtNJ5tHSZvd4BKyNPJY6fR83ncFsRoDGRyDZQdGS4pz1KcpjZnDJbeApSWhQBxStQboTy
RXXlrUVuSlp6nfmEl/yb8IfASBsT1GjqACDEQo+WmmJHLKQGiZxLW5BsIVv59P+UiLHckhEf+p1F
ZomEm0M9hk36Y0/5bMBmJyowUAZOjHT0KAwkZtY8mTRNuNRHUB03NxPK9n6wVLxcNSpMsqxkXs80
XhYwmux185iNeDjqsN/UsM5X/cK3KaV13L+TnPu/6snfclhuSx0M+7rRCxSKLFx9P9uQh+5DWq42
q1uunVCAajJXStrtZWzrv5+lvtQbt5/wEtdqptIHh1qoS53DUp9I7GjXMatR+MEURr8Q8s9z/abW
RDsVFQ9CJMw7pex7YD8V10/hCeV1P9m+1GDc45zqHTvGiy1G9ymNZfgWQqStgOWJVoDM8NsyR3xi
YW8+crY6NtDMUtRGs8hwWZKMZ2YRrGJk67svEean3ztiGdfJtWDhU/rx7XHqiorRFNnlQuhPzyKn
kgQwJFozbw2d+wuF/WIN2x0EGsZkgSjFkVNMCtKVjQizD41oAeSXI+GVE4VdK0fR8jqCf2FFHfwt
QAqW0rmHDhxODcmtugdqkoS687o2u+p/ADbLGt4/QFRq8nnaj30/IKgg3Aw1h8qnjkdlt359DdaG
gs5T/lI8F+l1/1JXzMG8ba/z45HlaNljKQvByJIBoKOtrEnt49uBnCI7SIaza3U/GFqtMmeVUd8p
1Wx9XJeH0uN7oJWq48mve2DXYJ4nALzSPg7qCgDYIheKj12o15s0DXoKD+IlcYo+xfcAupIDaFqv
7FFojbA0G+zAZwRuiZLX9/uHBsuTonbsm2pbxrHks/c9mJWuW309yRDQ9YUZaBxLM7ywmK9BI3yE
k3exZIYAa1Z1BwwtAbclwnBI0mTr+s0PnnSk0fj4xdB4fzh5S6FiOgNLyh8I7DusJNvt+jIyoiYx
sZRdkaVyokp8EPGWqpIBOEELx6cc9NhTrF+4uLV8oeEJ+mBalaMQ4t0wwtPGp+urHvG/Pq6Nv/Z8
cUTewCKXx8ADD1XNKM/dHvIF4xFkYNxVoMIwuNtyFLdZgNA+ABi/ZwIu9mEPh5+yAdupU36e3Ha+
+EonnfE6nt+e081wDYJqLQk2jeOsUXBKQZR4nJHgbg8pydxkK3Lrz3zwZ252GGYHVLWnIBevVWJy
WaDrpGpf46rRmCNeEFUnxFnEHMedxvDNrhmO7+2r1nan6+ZOfBczWflTgSKezF+XzksU0xM+SnYL
PlNe7rMingX738cPcariK2ZvOTVy2L1PQSFaMn6eocAURoG2pZ05hjZyOwu4JJDxW1u4BG219ajB
FMTSlfRf0OrNG4Jh5zcNZqg+rKZucw8DDBiUVvoQUoIM9yvwDuSPrMajnuyoJ3/uRa7Egt8UcoBn
FthjE4sXfGzubXjyxUWaQZ9RCNK7T5Z/h+ps8XtUD66ucPQSBfXiYMcJkJxYPKMbZHxf108Rcnh0
yGspi+CUCsJzW16NNnIA2kFLakWEd7BY4gUTV7ZAkw9V2et8J1fzVURkgoBVLweyV2Z8MnUImCS9
ctyIuLprLbI4jUwJFul8zGPerndZBFlvqt1KOMX04tplr0rSEbpH1FQunq/jQEZHJx+GAt19X/Z4
FMj42dMAKxtGtkiWFA6uCew56HmCaMLxGTUlt3vV22+v3yinv8VXtHa7ELioZU8EVrU9KOZAXD1F
xo3VsZVxtbp9IEkIKFpnz8Iy9B4fnsnssLWEyWwEPFj6/4X5OiMxZvDcd5CFG9Ks+Jo+9qDZ8Xfr
dUQr+tsa3B4Kt1/sUnSCRhOPgMnCsEN+ff+7W07J3LxFyphczGFXfXu1ohKUWU05eS0BpATHFL7p
2kByP1c1Nl8wvzoEXT09XUDdlpAPpictotLoIa7gvORO1hgZ/JBKCKpl7aQ6XNAuXngKlVUz05M/
UGPj7a0kXIgCyXYj64lPiLiY68w8NSagVNgo14zY3r9rASVFlDCD8Y+lrhrHl/4bQOnIYnWrnDO3
fgUHMrcLPb7asXhKRZTeGHtDoFxIvfv/GCTWrxV4EOHELgzlE3Z5gURNpjTzPMNztX44lNc4gSEe
GUm0AkqOtGoltc7/03PEjpjlD7Hi13B1QqB6efHJmJkCppl5qAGOmOESevk/UuM2zpdRTLwwNkru
Y+TGC2JoBU7UTxo/DTjGquudFncTXj758Dlo5De7k0yWSNJe1DB9wVvnoknrn3RZ6Qk8ZNwRAdmm
VJh3P7yTkpuoJI9NjS+MbBrgZFU3TEaoCwqsItjkShjme9sufNySuoq6QrQJuHCQC8C4aqAi8FBK
vO+Q4+CXy7l7FvPDJ3vCPPNNUuvMReg8DamEcFp+lweQyrUDmEC4lg5l5J4CNuWTjvGSFxHV5rMU
iuEZuA898+Zc6YSRN/KO3dM9dngEXGWUTE7d9FUs5T4abgrtbAHDfJDCexxz6brzYfK39OXuUnok
QWqoouKWHJAzYIj5sz3mRZOsOcc3X4WOFfLcTHSt31JsBEUlODb2MCXiKgzl4npbQPhwE0lQbnxV
bQeYb8OIvxYzCcRnLCynW25/fyv4fasXpJntA9wiaj0kBJwQIP8NmDfYoIeg9AUBHenRfJgPpZX9
tv0VvcjS9Nyb+It6TYqWzE+wz+T0ERwh/c/5hUeScSOPqgzyme4WP9+8WERW11vt3n3WNK1Fin3W
gS2AbwoNEzYTsQqJbxIwce8jmcv9ZyFovqvtOHBTB26koQdlvCA/UrxdoiAn1Uk+zlh8EXXwHM+Z
oh06smYU7W+tLUANZmqKnfW3mcKpo9H2HT/jKqLcgAZrx/tI5GpczNGzlmN2kqoFtsuwEM8/p2CT
vhOn6Ml3BJfJrw7/f604rYDHgAknU8g+s700c4BOEFVJWQJ05zrhtVAiaNlKRNwmgUr8TyxhIzET
UPL8CAQt42NnzuTgNDj4GfgQp/2bX+s5pEpj9U8TtcGLqvIFFFNEudte3uzKv4uLHFXqyvEH0hsD
ELwu8nwvjxhzd3A+2Gr9qrGbXcK5FXy6s6Bd/idS3skrxaDT0R30ueuEmJSNjmUrXpZBE2CRKiBG
6EmkDxJQmOg1gUlREvj7hFUaUa6/N7FIYsqLGVZ6NUfyuIQtM4sowRx1/IeSoukncuGI67xv2YzZ
RnntHLk7KcVzipa7aomO41Zk2fKAKl36PgypczIgzl2NTNX50tT6vF+CvFV90JS7WmEAOOHcaJh/
AgHLZCLjEhCPKPUaILfWJQGAmZp5Antpk9701cogAL/BRnUBNRkgNIsGxiEKO0IfbeY9kDP9eek5
Xiu5Zv9DZcwSotSJErwVSe+iR2LLjb/hMPR/lHfYykugYtouxxmQGp7bYlw1SstVEVUaj5xCcp4N
g72roIKNqdW3Bhl7TrjkHc/qYH13unNxTXUawt8e/ogck9qUaYTxe9KoHoO+jhrLcBpDBqtO4Eqo
q3CmQVDi90CN0TjZYkpJmsxHcl0rxp0SJiHZfhYiGM+M8A6NkhRWIMCTD7iD8iqow+2IhQV3Trg4
PCEG3dh3qNwx7PMW3bdhVFW7umjCFaCeZXNGVqzkGzaS4cBwivXcbrlFTGufh6N1OesOHObtkFZh
JhnwdWyONWtjvz2fMzujWFgubJhkgckmuXDTH8iDZokgf+bmLkDwSs7fRQhFoHtt6bxsUI90Y86P
GIXUpDO/yT/0rozV0IzeC8RUGNkMarIBHsIeLpl0DkzyqneYSQK0KXIWngZSqfTduSD2ZA+EX7lw
FAXhDCQH+5pam3oOfFFTOJ1ZNAO6GbuQHdSUpj0kAhxDwBAcVjo3V6H6Kt/7g66DEmvo6k8ygUPJ
LuoGe1i94ZEK6V8HaAt1IQQ7OeZZ+tKRG3k6Wq43ThaGmO4LMHL/x3KeBHK1tKql4jfw9sY33moU
WL33E3t4bnzUjw8r2ZZVLrROq/TEU1ewxIfe2PfN9ZDVxK4VuLgtWv3d/7ojc/lR+nwH+lfVqaS5
KpNtESyqGgWVc8yI1ArI9vPKmxhH1AWPy0ql4JkoAs6L4RHRDr6qDjJd5TWByQRxcTVCzdCeB46g
/7VBdGh3t1mjpqpjM0fvgoUuQW8adhQoTGuNRuFYXSQnCxJ8Ob0mZagnPj4GeGFRnWaLKNXg7pvk
DpxpT+vi6Rr34Hh30RiedmP4uEIIcPUYql9yFCHxX6nfrctUh/bwNZS8tg0qF1+HAVrW6NighLFZ
wLW9nqfyRMLup3d7N6QCXJajqVQ/RKnBN73FZyyQhoH5+i51U4LNffRVOFkUyDo/X1TNe68SRRLz
Nj27bbA91sQLKonGw1vS0/HUvtFLhiB7LxHI8GRXCh9qK1SwGAWuGf0gBAn8QF5/5AZahZSt4mLY
HEtwy3Ms79YvzuRcK9M0FM5W7CHsOZRY4LuK+dunvbKJCWZolusA2oEwk1BLSJLP89bung1DjG/v
ywAl6C4MJYUqLgaayFrq37ERSJFGlABWAS/W8kdYxFa0ii7gHEOzuWr+tcKUChakWuvoF0XqZa0C
QviMPaNZ8g0Vgu7Dj4Bl1zxlbJfeM3j1VS2AAc2TtbCk4UKXjNDRFYaDoK8VL393URugfuatXssB
dmHg8F71SiJVJIKV2S0Yr4p+DkIXLpP5WfSXSUbcSyygITZZYfzIZC+Q56RNFCgvBtEf1I+/j+NS
Ki5VLykqFhlyp/A1TvDpg2MRx37FO+qX6Q5PHanCZsjL4H9M1/f3G7AFsEwvoc1lWa9INji35hvD
zLzbnttrNEJtXUvLJ2bfZmBaDWn2EK4vM9XQPgY5vaXmRtPLqU1GnriEYxbINRq6fMNVUgrIA6gM
SHXUooYIZVxfGxR+0A9k3zK9EP91IqKjZcVLYGwW3rZDxWwY/xYojH72w+jwCGVm62+L62pQGZ1a
lNx+yFNiMZWRpplJtgBsRvsAywZVwgfh9d6gi2gwjgylfmAb4xPNyYKwl2BNppC0pZB5xYPeYjFy
Vuj7PxGEEU+NrDSgx54nVbwDHR/ERkqEjNEW+J8bUYX/3bdvuCWaLgxkOQZYRKOnGpghmFJ/6jwq
qXIqDZBvpUxMIDxSvzoL9hz7rNbPjyB7CsHR6U7IuqpzcPpeI+Z/BU6RfaUfXgLGBTppxLNM2NPr
rBJON5nXpIRjqNkVGoFD2WrptkLTu3iNJhGgrbFpBcKjuekYe/aHSbZeZUetsCtdRlThTZRSIgtB
UZCCPphpOi/SzWw+Ur9X8M0+dM4ihsfJwsnbKXSy9+D6nXQihhLexzYxWWLkdIgOIGmbHHs/1rrQ
4AzlOcNV8BKhtPXCqnXSGG5JpHyAO+V7r+6W4fomJ8flim+8Yz7YWfAfeqbm0QyhQIPXJVVgJOMr
QJdoxB4Ga5CNgyXR2G1V01MsACevNid0D1xKruzZt+ApWY7G2X6vjDMwzLUKSPWYg78SQ5tL571r
ObG4SooCeQh6V6VUTbxHRJWSvce0l4jtRtknBT2rxZfkJ6/c4GD8Q6flrdfXSX/Y9peFMY2Rv84l
NflSmwW/T18vP0GvgAx58+dba/bI7xQCJG0GwEafkrr7tCs6aR6Tuou+CxkJEioPuXGIkYksHxZ7
l/C33slOfxDF2XP/Vantzylkd4HtSRhZ6U5NaLvqGvm9TIWVXwYMUIe17TXT+3BKRX4cSqxGQgB0
dJIKGgCsFyxt9RWKgMQaAqVQh9cd0GIUMS9JSA4E7diluI2r/ku71fhcdGzcjHWDfQXReY2oDOlB
TkFQrW+TmoUpMomM4SRVeAveCxeJlxfrLDUQiMyKoWDOBLpqoLcUAP8xNKwGiFjw4hFYhF/FpwUw
8rwekqwZ3LQJPy35tNnyZVCCnO5UxnDE+/YMHDh49HY/idCqTEETV8Q/f7pRWOURtMl1FZrrO1+v
S0YI7UTLGHdmWFm90Vz0zoLOyRxdHHrp3oL9cREtec0ETdAGz/GP9cYxBmZ84WKXMp2mqczxKx9Y
En6SirDLwxazVa+EIZzoth2X83Zl3of59++Q0ZR2mOEptt8WIOgPTN1NvTs5yGrlqBXXb68Ofrmq
RMhtNrYRd5Nxl0N6mwvGz277T38+Lzurut8MRfKn3jZMrfT6qmYpaQo+W48+xQ7Ib1ZlzLgvkh60
2fMlFK7U6RHdRjHFR34JXqxtKZiDgQZlGSIF0oAiVRcnHbMNOgFNdozFyoNaAILKL2VVaHDjVyV2
ZC1OL3MXek1aV5jV7UbxIXzHZGBQ5cj+Dr3xvonvpw0ck/3QS4Onp/J6QlKdU166FgCOzM1OMbFp
w0t7Vcw9MIVxkapLZ15nJ4nkiNUzgUrMNR46JxyX1zxn5j9T7un/rse1PwuCFnEAaIMbb0Kyd6xy
LyOxWfjP9wCzwfZf9X1Iaoes1KYzt9rWPBw32rs1lh7qpMRECyIHc9ZcKS7o4DnNUW4Mo776MZzE
lqrLwI0I3qHxCm9Q6WknPipEJpb6vUXQAwVIg1fC7jup5Pb5a7coNU8GgbftvZC3ojS/crjJQnNY
eWxSdqLPXZCOJrBN6W0/eU2kXPfj3+ueOs+lo1MhM1GKSxTLci9dODJ3IhR7xPO/xg+DZFB3HDhb
8Nhc1gOCiYM+0gTB9DKYRWEvvJV0JkvMxKRBxKMzBr+Rjjdi27UW1n/9mybGWvHKoM6Fl7znYZzs
bda1NzT75HOT33dKh6QYRxio+hO+ekhFSf7mEPJt1MRZTFGNTeO8EmcJWi34XQV1RdQqwBAQqnPg
bUXzPHcMCIInXP00F37cj0WU4uZyn6p9OxlFPmIzzK0F9bHtjbUr02G7dzTeShBPR5O/qEtH29FY
MwWVfR62B4o0bI1pOkNY703xFpFM4MXbnG9dh6QssXHLi4umzA8898RUn8u5PPHPFXdkmM98ivz+
cdi0a+cLr9S5a4f0MZkbTCtXgN5SKddbixXnmB8nb01JGmXuydgtMpAh3t4dnSIPnMEnGjTt87j4
i3z8VxJhSb39w4S67cudDnFP1EhQMWY6oRrVKi2FlM48M+UUQFv5q/qOxtE5AdNx0EQidw2KU3x1
1JFqG8al0TA3sXMOFg1C9r12BU9i2syXQdu/YcTMj2VkjLJzEPY1wCRQOn9lv3FFGvfXoEXr0Mhu
BKQfsj4zdrcbo/X+sYewIWPN5yqKEYu1EjcEY2qoyOy10UbGo0u24/Ec6x8Qj+3ONebEPiAugi1H
d+/eDmWavMi7SfkJXD81JDMk6qnPCaHTerCv/KV0ymC/MZhJXepbLaW8U+Hr/Sz3ntjO7hnCuW5L
XF06Oi7PhdTOjbpK3GOKdAptf2Lm2efmoeOwUZI2GHdL6c0jJC5LsNtUcRp+JLZrsdUti4GW4x/x
W2E5HUwcWkyE6YHGH0xrGbbR3aJNYPz3vhAMaPJllmxLYf7U46tLGEguFyO/yfVzagAip2kIxq8p
FLjXWUqjC4h3wpFPBe7lVcRrSevfIl2nP+/yG0o+sDEWr+Q2hxUqQB0qPaXfIkPb4CW46DFu97vZ
FTBU1fXJZWGlkIVACDrybJYCkcafm3qBnxFvbCq+s/958apigfsiEAFjOPqwz9KqYMmUkSBqpHxD
hbWSyzvQTDkcQFZmYQ2yMZVVztkJnHmJ+pWkD3cnCzRQ8bU4npNQLcVIf7tcE1VKJsiRhH6yyvv5
9pPuQz0yWG6KFcVorDfp2GhMjOo09FpSxvn6FWYAHHQR1HXcip2HjysHh/4o0oLCoSWIAaJPTN6t
mrg/X656jtKZfOI/BX9DJijIC5wUzz9l3VidImzUJpHUoKm6hCq1DGCDCzmbwYxMyOgPL8QTsAIL
etSb6OvAZImNiVbVrVQSUr8fV1ruB8eIH4+4TvjAs60a6PjKL3ekB4WdMlhMG60joHYGkXWoO3IB
E3ZB8nsWbkZuQqCLtdQynL36WkJNk9g2sfMrTUSu9AMgWA2Kc2ROpOiJ+5neLtC6v7JHvS3vyobQ
1+Nlqz1K8+A8VtozBf09ZSfIELeIoCUqgzSE09zSbIifhw7EHltiHMZqqMZsSUmcN7YAJOO5dqM2
beM9ftXbLnaeaCneBiwSYIOcPyn1aWHFoFiMMndDGJVQGR+958zK1QWGDUZyQq2UVfKHwN0gFORm
6/Oy7p+iwr6SEZWdTzB4BwCLT09z+TlqKAHpmt8sOOmup38yGmYqQl67WKfej6CGfoHMPfWGdR1W
sjSVe9ix0gcAIGxTkW6+DC+yYpJUvx17Rr0WjnDZPEJ2gl3bC+sWu8UIr/FbMxBhqKfzEQxudnDY
x0Ds3XEHDGwlNTY2UKw4O6r5i9oiV8SKG3sJFbx4F7jbOSJNIcjaUODCmH+q7V+iU++j0zEl3Tnr
+l2OoPtjf69OD2CZuyeYbL2duB/oElfloXhopyI+RSPLHxVIPuQb9t78KVkG9SXUyBFBxpoLJhrs
qVrAzKp8hUFsHe2CJqhZkDMO0+xmX44SVhWsO4ANsoyyjyfshDkp0I4D8wT2PC75oJK0AKog4S/X
2IA1cA+vmgOiG0MN4uPBHkZRueBKtrz/aEkkEGKssvklmP/RThqcG0SuaIGD/dTjy2QR2okkT2WC
3E40MFoLcbs4rxlVeNhV6Xj2XBws/3xRbaaYdtJjiEoFOfeQlHnjWELpb6FgV5kLIommzyQfMRLO
jWfLZbPvpxO1hCMIiCWzdHws+tqi8O2xTKzp2ElJ/yiirpVImJWjOMbTz39lpv+dJbyqQQxBOr/g
VeaHlAsMFSNOp5emIg42qFEwPZ5JHm9AZMpZHo6jl1DRl2eE0rrvSuR/Kq1DmVu8Mib/m7LqmYRC
Q5oRLUCxS5hh3X9JsU2tF5RYnsa128TKOlFifDzECpuccyLSK3RJfq8/4heFRRiCHHCHY60h87DL
xbSu1KxktRbZWWprdKRZ3RL6y23ItVsicrsI2Wf912r2q2yZ0N23mi8o9710WNMZCnhsYr3g6Y6w
ldWIEavUVowEuA6/CjbmxDg9EZIQCKBY5yh8dJzT0VAahVPm4KgDYJy6sgI2rwUJ1DUtNw6z4EhR
lPyiFAX7C5xeMEnvteLSoLJXyaaszyCNTDI/w/LFAHknA+sOtYDNwLumQLeRyRW3Z89CPRyPocSk
8QG65QMvoUhC5vXp/8+J1V86Stys8pdZASyRHXNK6SxPR7dwQ/DSqD4mo0t1JJZ4pEa0t6KlCisS
xn9kfB95vcVXOklii2kpKEInlrAg8EQlDIpCNdzw7mLT6+BGtubPeTeJZWHtWwUiTMSaus/3bxv4
Etel8yuwzvHfwerRcSwXzWrTybIHxXG7mCORmmlYoPIcvVsroWUEbn/erBuGJL0rJ4PqeNVcwOTO
yKdZNIdTr9I+GdpldAkvT8PdDzM3KR7BMANEVH0vB/qBZklQEaO7xo3puQv4fEbaMPMwohOCLaHz
OYw8FyUL2qdCyKabz4M709X6uAMhPRnZ6U2sV/M4m+7fjcwfNKTbZyeckkf7Qzb9YWn6VlF5pVqJ
ZIFKvzSXwmIVkIVb8YxU5tNm91VITcL2XSlsM0vYlsn5PtJ8t1TrLYytVfwugX9bHhzuHaWxwvJP
ZWhR6H8exkFSgzRrBOpfIO3YO3LmpVgvATXpHoU0uqsPYwKJtkDkdrUcMtGR6/bWgHl1H6Ko4HH/
9PYn2c6cJS3mHPZhAqvQn5srO8WDxQiNpOVQLxNYi2lOxVLkf1DD1DFtrVa2bUT93Y/bz4Z+afQs
9trTR9OwRZhRfbW5ZDJjTYAVSHN+1zq0ENLxKvOqOJ3uWhqzOuLF56eVuTwXf3rROtL1UQTM7OTL
JYt62x5Cv/8yLhFrmwT7vdv9U0HgTok5BaM4LoAU4m5/vL9lKCdFWyF+nDo3i+nEnjCjxA7k6g+y
8Jqf+r6KvpHkgnjef6QnMUgo3CGUruteWkOmymtSK1jR4Ep7gAtDeWKEHvUWHZ8Y7MH3z/D6mTcV
FsfAFE6Tmrmeny5XckCl6zO1Kasz4SJ1FMeUOcvginxB5/1taFGquCf5rvIYBQ0M9ajAQ+01fUv+
wKhD/cbmpOVseiLPq3KPaMahYcVbFHWoqCWc6KN/o2zWFq0RSlQSdgzSwMdnBFfvjzIiHUmOIl4E
QAnCeBPsC81P4ivZzPJ8su9qCF3b9v5f2WQjyU0Hvn+7Z3DG7M7mTtT5NyTXzPXk/BzwKG2BW8xV
7WQG80wxD0ytNiI5X9XBaS9FVVlbu1cSCbNTfJeLWHF2RbBAEIpwDNTifHXqFiuYKtXt9GjU3pRj
iyh18A7EzJADwgFFVtnHvUPan8cqDJlgcjxzNh0C5or6CMDtqGHH6nDmGeh6TsPVTv03G7wa4JH7
jkRTth+b3bROwggkk9WSherciLLL4KR7IBetirsDTziK+by6p86UvKDSbeg1TBpQvwBIGdhH2bkT
WWsokxJPfCdNqZ2baIBX2Yl511ea6a0mLznAr6EKvJZCTOTKlqds+GYjfVUdb5tGjeUTdxtpsoYy
nyo0WmncWSjxdLzxtsveoXiRPZM8oA221LO08BOD0/aWldR3nxsR3Y1/TO1hoC7sSYcrs4ShuI9B
Q9MHJIFLRdhYEa5M4sdlmkOCRszyDaETfym1OdaDlXApfTGxP3bqDLYbiCGvkyNtD3estf+sfsCG
mqtSUDQu5hKlRV7KkpOSu80xOYoKFQmOrvh/EfdItsx5Myj3ytiCtSBBc8Z+aeQ/qrePep9UGOBd
B+rlwmCpE6E4SYVsOWpjdkLKRkdHEw3LSO1uqWq5I8cSryQtLf+t2JGu+6o7nQhRStMqr22eiTh7
rVo8LL9Nq/6rTGUUYkbmdoyg/V2r4bwzN123Md7KUPGUJm1jglFNtmoueqr1nuneFCXhEyejWKlv
FFjUnxbQXhDebQMsn2jfnNJ7q0mNG292Fdf6uhplL4jiCG8AXJoeh2YUPCmAB2OiuOjUTHgRzQbS
zId93XIn+VPEF0p94/bOR72p0lSJlYjbplbmregSdSqyfwOow5mJVsIK9YNflaWPoIhyCwwMIsmA
iCmJiQ/lJ3AfxFyQKUE5L/sIFdjzwd1aHos6XLqjTliw2Z4CsG1jehvlXmb8CFH23SGNzDOqSFhh
uLD3GDbsY92y5L63HAx1wkpGjLNRaYLqr90dT+LV9HKEKpZ89Ho5Ce/xF5ijkS5UrWIpfF2dgTxS
cW88TZhcZLkVVQiGyMkpIEPC6kUcaEJVKhcc67N1oHGaslpp0ODxolrUbSPc6WiTDj2BUv1bhjMT
2Y8kAnI0B9hpBOXV4Xo4R1Njp6ODz+zPldtrg9tqiduI489lc5cGvpJiQCrKHEVQ0T/LDYrgEP+/
WqBTCJwELdvxHkydyV2QVBy5LumrvHDcwn77dPN8YML/QbzqVpZfcUx8P6qRZ98Ix0bwIt8u/4Zv
0Svlgfk4r21hOyDrTRcQmucXPakyYDDZG+YOsRHN76wfG9ZNmfOz86QpwjCcy79wMNt6NadNvoro
cBG7K3U5x+G4PY3MCbUlDtCc8g8b/H+GciH3TmN63wksWNlsNKD9GQ8K+NokI2ZO/akjFkFIYJD3
h8itVOSUpEMkC2jyi9jGD5Y3wUE+3EAC+WuUha6pdCmDC/Mjb5YSA4p6sMPDAEoRnXKmFm7VUBal
fzJV6CawexFc2IdAjChxNkG+yGolmhiTb1rvdCltuQi/jJwi5U0K+wcXzhw6AqF8p65u1Mz3YNqV
k1TZC7ACRi4mUf2eu/Q2zYuRs+uY6JV92oZ+ZwaLxxnfntSHcpCt9LDUHlcFtpkfysOd/PrRugCj
ldSNA2LJNk9EkGv2vDv/RTzODzyyPJmn9+QAYvxl/2XWvQZTqFwGqYaasoTnWXAS93bCT6lgfjZs
4LW8zKDKZ5BbL7Zb1bLmjwDIDJP8WBKXdwR2YiNUantWq7uapKiegLbA/qiWUqJhBM9NQgFwWNfm
cIXGYdCnT19kauetOh5NvrBsL2R1FlNxgCGiMZ5gRfbaQTC7es8mhnvbYIcy8zgpFwfr1c7xBzFV
2ePzb9hZLGlySXIx34pz8XHRV8sVBfW8sPnnKKdowGLmo6HjTjBXaz9aiT18/gV6BdO4VredlZUE
rJs58SnW8tToDGHzIdThsUgao4rUIo5M12AQkzlN6xGyGmjRFul8g+lF4boVZWjoaOlh5g6oXlgk
v9bDwhNWB202TxkC9gHi+3eCdmqOwsl0LM1t8hHzliL6kWBlHpcRbLGWzzeKYf0U6V190OEwjxne
RHBw7dku7NbJj+3gdEpxycAlBGzEhQymfw0BnfkAAWN9Y4vFzYCO+Du+D5qPnypvTAOCRumNFBMh
+XQ+WmkznFl4rsqaUbsIKYeBOaB07FkLfLz4UiAcQfA88VUo36ay+RZdpZ6vqSZ7H7jDSA4NbxKF
wUQejNQqRp/rnoyuJE0cBUd5e+9L1cdvrZ9hWcBwaU1eraruA/4PRUADrMkv2+t8bwDHrWxib9EI
Ud6b/EC3STljRey6oLQYsM9f+RTDHV9zixJ25Kh0F2W95ZZ9aVSqnLWof71QyVtgCUg8pFU5Hoj1
VScw25a1QfK+2syA60KrUSyqGiDfyxQ93lx10wV5VauPlaB+U3zR7CaZa+XU0QZRisFGY6JfI5cW
2tv1Vlq2rGl0QmeM9LiDZMkqyzMXWMPz0znogDll5P/fuWsyGyr6L3bAHAGKCHKsWD5ba9cundWo
jlwiymj4Um3mmGDc2ExfVZ6tBYN7cZfCYv/oaJn5ajWFvCNEwx7jKI9gHmiDvSKPA8CWbOxcVST3
0e4MymqHjhfC9gZ9HZLcKx2y0OnvzX1RdccUXbLgtw471ykSU0nTINJr1jYelncH1ONl4blunvE2
RN1efiuwv/WqnESgq0Lub87YfnyYIbZcnHfzKTqYFcRjYCYKK+a3P6HawpdBWiDYYs9WQOIyKbD/
as3S0LHDfbbuqm88VEz4pfyDq7dRd/t/UptWeF1TYHF37fR3YiU712mija9ocj9C7Co5wrTu7m74
8BqfYjzMgGPevL7UpRRbhttlE5gHA+NUbHP9PqkHfljKtQv7TBcswSAtpgOZGJbGsJqPnLOJDCPr
l+id2Cqhppsrhj/tA9HVsr6kgsxGJpwcJ7tSfJtwnCkZwu+urUsVU5HGOBamUxlTAL2MpQmlpq+P
AL5kdUpTglEv89mdUR9+VJpUNdojdWfNkziIG/zEral16j2EX+DFcgRp61R2MoGjoG8eN01R+d/C
CsySnvsVeKM2e+Z2jSM3/49OTocTC4RlPFB+FMuTqz199ZVnDv5RmS4qmnKdzjKHYKXRfz5KqPyG
g9cLp6r91Y6D79Zvi711FPXLbF23ujvzsFUSRvurmAFcglm9MX3taD+j7WewFmJ679QM1nha7J/V
6zj+kZoHRthKQVUr6eZkobanhNkcCtkqu+dKHNDeIl32ixQMBjwj1hJ587IyWTISr5j52+UibLwP
OS9p+kaX1EMANUAf0YqW/oDMhb9Tk/157XwlQm0G1+NGvAEVmv1PYGiDo3Ew6bDhE4ukvqfl81fw
VNsfBrq83Wl0sO/vH4FnWIoTqPMTGFeSJNxcGvNXdrOs75zU2RY2heKj+hA+igB0scBb915xAKzX
AgRuxU+SydSh1lDFTXR3+6utrYSjOlfGolNPcfBY5Lx/B13UwD8bbrcOlNLTmIGh4BT1TGJHOpPV
FIK04aNrYBS961CJv9UnpA4+Lkt8d3/aZ8Zt6r+MoXTAp/biRBwPL3CMErWva5Q8hgSUjdK6XNYO
0Cg1onn4vaZp3N/Ap9ZoISNO4G/LRAOZTEZP0/GLkP+q494oiG3LalTDn7JM+LMn//KT0O3di0M5
wYKQqz7WBpKprkMDu/3zNMkS4ZCfQPIbvxYkJyGE6dZA+1PU1/Glbvbb9RPRHARfSftgis/sYeNl
58Bb5VXBjcxHpG24FKc5VEvOhlqjsBEN3Ikv8dmo/0WS50VxwJ+1hxsesSy/qJH3XSOtxDNIxPSz
QhogqJsZXD4BGb+V3IkWf2BXn0qXTEx4NbIJUl0Y4EQxxWV/EKK/deDuExek/ffuds0qg6znBqu4
gWVUZMaJANLjxu8PmlEfgSgoPJ9350vH8B7eOgjRNdC8ws2Di5NF43+XHZ8iEEcUKuSutDpqcDmn
kTqHe1TYKO/x6+MHRW5c+WtxxDdSDdrF+GrXqQ0BjiCPtBgSUwzWfQxi0xdSQpz1iai+lYoNe/ro
560BZK6y7LA9+2ZNB5VpuTmtolDA/nX5zCPI/i3CQ42a0MoZgJy1LLIPSz/ABFT7BooWUJK5V0OS
yvv2a4+HIWgncFWmNhdC9AaeN7N0Qk4GQIG6iUYWQHuGSQWHBAxh+Tswuu122g7XaqMc0jtI/5NJ
YwJuCE/1zBI4fjZsu6vasJSV1LutkhZ2EQAEwnRfSRLl/iWgDhoW6rMpOzrmJkMsoJWT8QjwSA/9
h/KqoajUzcXacbj94ADLTG3/S7cwR/QNv46a5YThU6ql79iOqpgFX0Xqarq7AO6TnJpa9v2PdTLH
IYSZNSQRDuACs7vtuUfTrvcFsC0I8QaLSMyGI7cVFxhP4vPLprGGqCJAp0AVt832QwJfGv35s0cl
ZKaqdjiNXDB5JGjR+cSFO/mTaU33Se7dOCCNmMn2TM+mrHImx5903iI/i/1s13oUHz5ekY9umzlZ
I2FCEz/79uFCIgBo6SAu2vx5QeFU4TAi/vf3KTAbw1g97ybl37g+L+YYB+NM0wqg8Z3X8SitSl99
OjWKU5vdRM4xjqk1i/DtdFO/huiHC4BRJ4Vyxh5k9VIsAmCA17/CzBVeY+WjPLcTDbNNNCVJf5iU
tH+pnShT4pUkwUBzvG9fmkzGcZ/MfouhIpNjZJdzZmIj45007JO0mp24Odr8Fy4iJoqDtf8OEGcF
BLoxxmzSJqfGqP1rdjrXf5kJ6J9H9KSRnfJwFO3c65XgozsnNLUOclh/GbsqtpW806RS147VZQvb
trNRAnotIYyYXcIdKqScquC7mzCMztYNh/w5bBFmeBF1dasyLxljxu4gp+r3KXAwdOMIunRYfcsf
SH0zRDj3vKUbez/o/LCXDpFWTgIMxuTn26AttbiO0S4fZuiH0etm6R30UPw2isv92lVVx3YYjR5B
b5YB8O7TN+/vep2Aa6qTIxeLd4loYIMwWhLVMVvSqLZ+72tjxz0chVzwqkYAtLpaQ1gqn0imneZd
XNqpbA32yDARTQFqSPyDVsMf8CUeiA/fh/HPSCYZFNj67mt+XM4DvnFVQlfvcL2OWfZjdSlWHHp4
6CJZSSLbu5XUp0PXojlubiLwT1sHJOsTNcI3uhq+KbNP+egaWyucl7K23tiorYXwGwnHzfqAiWJL
snZ9LNhti9KeOW3VSQpSU8xHdy6w7O3wCjAkhT8ZM8oWau/GtFtIEjDLmYAicQr8SZRL9kTxKs4F
AAQUdi8H238D6i76Vr18ZLuj72+bd5gb9GiSeUq/pVxWyp0VoJULpqVy/EOWeV9xGLmrqsAXPSFO
hMWG4+bunafvbUMRT5t3t1HPDkjHChSLQRn3RniuMEqbwhH6DSjesRQgJLZD7e8yLzEBkaCtfLqK
MdFcb07FguNiLrZN9XuhoWoHD6AnVT2HmvntgHbJ6i02vfqbV3khLH3ucxaWcfaz80gEbNWWpFgt
36nKUgDBMCbCW0vUL+hszBr57kAgEI+WWza1dgQCmF7yoGmXRokcgQGneJPrSuwSUXu1V3ZCMAMG
Lbsear0nT4B1kxfYcD3Ri4z1Uws4ZX4HYt2JuDzCbtLzJHn5YnDEiUyv6d57PwI7Rf1LEfkJX7oZ
Cab96+oKFm8wFBiuwmBXc/RXTUUt9TSvlUuCI+FOsWxp7pbEOdnqKJuK7eoE1u5QZvQI92d7odxf
CtC6Vw1Y2uLCqQVNehy/FQZ2XpcTEkXebiQXtkLLexz+DfqLgbqCHFPjqwjtIN8re7nWeaScyX51
l94ZpsNX+AHpnyANlPedYw5fsxRcT+o2kSwoU3NmUj8nP6T3LJ97T9QGO2U+r9XdU35ltBy7XPaU
FpRSiWXjSF4JE+bqx+Nhxio1yD8qgFGacRg+MZIJmkFxwkpstPQTZzso3kTmbbFUY8iEzc5M3d7a
RMRirAKJ4TuAH8lCHZM02j7H6gpmb/mcF/3GKY2M4RYoTaOP+VeONWMi1miu/diRPjPOwN25KSBI
ZpaSJ7aUf/RdP5h3OzO9ysRYfMSr8wOdd4Cj8sJ4DyGCnHhjMkzWfZK3GGufkrd7KAcVXGwpgkHv
Dv1WXPvCox7qd/ilsHDcpcpYXT+bjMmspdA5s84Tp/h+djf8vhdbPV8k3vidVkapr+1lEG9ljZsi
DBcEtevpH08yX963JK4BKJ8r59K61IuAlk2MQLMYAvjh+5U67RQXX2YZ5VxlXdDP+7leV4ebi+4y
HDMJ9wgL+JcszJPzPgnRzZEdrRXB1xorXWcN3iRuNM3P+cCVPniK11ZEGwdr8rWOMh3q70lK/F1B
3aRunZ0yRVv4pbk0hyPiFXbD97ZnS/bdP0MgmXbyk5jfK41VOf59CVgDmeAnCj96CcXjuLoa6A8b
OZa+L50Tdrf1A1i3xa9dEnXgJVaD9k1s0GBx1M7gZMZ7DKWoOe0zVV9T8kZAGCWF8Syvsw9mXS3d
ziCM0LE8VI2iVwDVohZgE0//sr8lebIgqgztWFVP+KJq8xLfteLIs4Pqb8pBg9L6w3wrEq8p/B5s
npHRtEIKefNBn3yCRdTSdI74SOx3ZJyIRPQW08uOaPq45BIym8symsy7zWhsSpgquDir9hv+8bqp
xoUcxQQ2+kHysc9K72i1rIP6bfqAvknEbIHiBe6yK8GGri/BXWJ83H+CbHv9YBKPxIUTg/YMbzPV
lYA0hBFxa0/dahMbfrhn9a4KMJ04VCrUjqQhnOoZQl+AvKeqNfwYJ6oYvqZuOkAStK+twsLcZttt
ySLaw2IHPeEQuR/oQD5eX50mIFVH6w4JtDxcKHEeW7qfl4rPezYKcby2+OfnGSk1M5waLRMjKl0p
bABRmC7WFG3T4cKRI27l99gx69Kzj1EkQ3J0M95JJIpqRHyW37PSa7/EVca1rNzNwsOE6k3AhKdX
5P6v6oy9yXOf/o4OadsE/Vqe2UwByUNn3tUrWVboD3xhFa/vfL959kJ0h75agfYRX7uNoTRL+WWH
clZmMrtbL8oKPHYagNXgrlT1XyE14ISaBjoDxd8wOsxCz4gSCnTscsWFi+dFYlvvmUgfd38cqqF6
+vI9gL51dOwwQwnN2O6reUhA+a5XEKMelXsxoDHMIfwZtRZPBDQXkh0kQTXBhlC5MPXAs3HHySi3
crayWOll6l1OmixTsgyfstjl51K081E3nXjbcaOHXwmQRdSz/A+wjgJuDfcFgQ7KTf9H5nS1nlxR
pGegGdWrtvyMxjPX2AGcPI3+s8dV2OGuM8dNZnXKYhnl43ea0kM3hL6MwLiaEHahpD32Xx6ImWDT
v65cIbPrvGsCdFJhfgpjXrGxZTAD0DajiO0DR8SJbkCsOS4P9w3besY4Dq6rqNhEgOZXqxXzyqdR
dbn7zWSZp22YpSXA7UG0h7BA0Rh73N5vz5SvgKCutPgQQrZVg6MKakuWVYaH5pYhgVQ0Mi57QoL6
vvTGXt1TqwlvNhW8V0QbTU3Oya8SMSKjPO2+jmJgqz9yb+hzASwD7I6ikhuOfpNi6O0AZvzMtJpx
ce06dGTAV2Tlax4kGD8l3MzZbmlx3V/i4pIQKYBgK9eE++2gyfAwtdTDIIwJp61NslBiQIYmeIC/
NSJ+v+P2lYitzs8hLz8ySGdfzz3ldKJEvXZGpdzEwWSa/mqS02fGSXloTaI9DSKfpWELJb/zvxzF
X0hQ3j2/S0Aiu3bVty8VTmS3VQmx9ULIhStZFpmDbGCzZqVG2bz2I9DlaVtfA2/UvNanJG2bfCnt
NtNYwp0dDV4IXjzNbyveImfLMBVlwQ/Ym0au4f6LOU+Ameuc8FpQg7bbtZ6AXNagLUIu8dp+8FkX
+JU1yemNcrZKazjzS2l4Hl2c09r3aTy7hfvYhmD1EUEktFa549GXkKS3zh03GE+6oIOh6Oxr0uO7
bmspx9Ejx+33g/UN+9fffGGiPYldAw7i10zx5R9dF6iiZKVKnPFoLnKgE8EGAxT04UJCEcstOZVX
2a58z9R2JjKNfS1fGGGD7TU8IfAWwEzas/WozH21KgTLcv2QjTSquAE9cSKZBK5KMDBmTIcvgfln
W1SqR80oT1CPIRO+qVPJ4qAv9SOSR4+SFpRxlRaGHRt3Y1DG/do8mXo4bzNWdA6RCObq1AIRMLPK
vgCmp1fkKCDRmOqaVdlnEV/LE6Nimwt1MrzJ0I6ir0r+0gtf8Ds5DLyiTrhz6YppZp5unCLN+VYf
Ko2RGHe6L9BfhZdSEwVER8Z07s6illr35veNfCN1/Yk5xwwgdb51CvfCi5wW4TrG8ScZwn7ZV+Qa
PPebEiyaJFvfhoJg3o1dgfIyRf/FvWNXCKP3hFfugE5eI5Kyjo2XJodoop+GOWKSiFjnFBlxUqn2
JgtICvZWud+gqbNHzdMCWwAA7kvMjKNdBATIXwbb+4BFt1fvtPwHNtnEUKz+XewxA91q/Ud649Da
8rtYjwMLD7HZM2FN7XsVY+2NWiGsNSj2+GUaMzAhLp04EnbvXImwSUlzgdRXRKm5MPD+Hjnblfea
+0yI2ZxepREnKF3lUKkN2oBwp/Fnnwd+xS/NZlKHbabq15a2qkCO9QKfdgFWf7Jz45GzdFjj1dq7
VCuNC0jKuEa3J9ZApwB08B9yHWdSqYbREfDIQfB7jddR3j4HLWMPci2gZuW4HpD6E4rtCb8mBZf7
kwSCVcGMLt+gPg2QV74qxn81zWAZ7IF0Oe54fYF2Y6/NAzFlfi0gPsk2zLrPTcPnEPxIkyFdwjsG
ctWGWX8CV+q9HGTen3XkH6+p3fQsjrgtou+2Uw1UrVq+KPuoVHhlctBJwmC5wlZ4+gahCKMRSxx9
fQ2LUrIAbqOiS8+xQqXIGsNtM6IPztG0aVTwDg7exuEj+Ow87xpXiS63lMNfdenA49a26ClWAuR5
B6OzPqjB1t59lsKnRDyhemwP4dMMrGPGGzpWf9yRRZ+gGPDzC2CNnAOlwzW054RyuRh1JUheqtxR
/M2gIH285O69AzVm1cWlmzN7/JYeAVFNfHyUXmUyDPkKBipkXjyu4mBnxVL8mZqVBXeHGgwDqP33
pLL+g9cglZDohKkt82VJPPN90hGB63e3GavKIm6i4BgvqiDjMgLea5q5Ig/Kzlew+g9jonPbv3VB
avSfy8edilyi+rx6Y5P53ROpnVTyAe0hdpqHc9H6HlaQR4buk7eAs2yOYQGpATCXh+DPiXeQVqeZ
dE2sto8rmx605bMW2iQ3Cbp3lCh72L3LcTC88jNGMGgvUYITpTKPTLrVcNaEER4kVrtvAA4206JG
zxCKGIDASgQ0bvziOxGo9A4JaXxL+6yscEmi3dVjAYIjhdxtuOKk3oAbzXpEXvQmU/QiNCCUqeUQ
A0dZNrd+MC3MvEetOCULuWl5C3/0uqjphuXj7O9RpxAxeoxi+uzzsy837oPjfRYGn2rtLUpUR0dL
Dh5aJPn/oYCGYzsBr7EACol1TS5pAf7nyxfaz20YiUW7qRMXSsjatizQhrhoVfEx592gcA/CxJhc
5wHFdBMw/rxJj9hTD3nArNSDKQpty4GmyBa7hih4nR4DtKq+dh6tG54AgL6jDpSrX74Z811OaW9/
T0orrgqjj20f+VsgavWOjE6OnjJB3GA5d2e/Oq3SQZRkkGcm3J9OYCfdQG4ufihizscB0z4fU8GR
DicP+/jqakG5wNO9hbmnG1iUppELFH/Lu7SPv+yTpXhN0b+6m4IiEypqa8Buh9MM43r/3tIAlwOp
5Bl9XWFmX/uX9ySQmLWDvoByTWfTC3su9IEzfiLIUlhfs7tj/88U5QBn1qyUDoBmQFw5lbqqSj+G
nPZ/piheOhUvdBDiZn5EvjzywOIWe09S+IwIat89bPzPR7ldScm33kDbcI3quR4v2yLOxJPVFAKl
+VRQgInYSYnRC4isGeiTymNLRiQ/F2neYoxc5JNjdxz8ogBj8R2KrgbsGn+WnmUsL5uAh0N4jMYa
Hvy5Jab6+BvL9eoQpuYCkc/yotNA/YM7p9hRyDnLDPnUw2dDozXblqaFHSmSoTReFWzviPmBQshf
XqKYdRy9B31DslELfZLDOeQ1u4HOgtaUPy+7Wi5jdLPwSTQlwqsH+m7ki9iE+RrxCbIic9bnJQsg
diP+S/53uAucOnu0HLShLXydJuEU9ZSacj6ZMKSO5+OskFU06iPL40DqQO+YIpvDQZXVMeP/Evcf
NXCZdEBD92jpG1Hl4+B5syqW1fJJSHPWR73EoDYnKnDc2k1LAYatEoC04DDzBde60khXeqpGPm9l
0sn4EhbqLNOxCgMibq3mFI325ziLmbXvefjIF1BbR/bivjSSGq1r6kAR+uflitW4x6UCfM+HN8Gp
fAIFh8MULyeetZ+EBDQlXpdwl4SNOdpYAHUTlZ9hT5AJQpweKFsw83tdBRNBTV1GXLUsjjtoJfPf
+oupajGoijQoCBPHC8MwcGeAFLA41T4740/oCY+TcD958Zi4BYGeF+75QsdcDF5bHSh8p+H0M4l3
C5y+1fTCz5iHTwzW2HV3yk/XfkgElcRGPIFuHB39fNCvSS4Etelkg1+npKbXH6V7gC68X8Zg0rHM
0qfXR4pELhLompGQumkuAdX2B0MfudFZxW2pPdvMHlTGXcUImjXrm3CkiAdUUs9lp00Rvy4OxXo1
DYZLVeZURz0nQ7AFPtuCM+4+1Yn1FcH/wTObDFlDEe2+0i8iu4bZ7PkxvebamF4s55qHf92+p/89
OirzUrdeviMnhwBX+PMfljzxcszh/IckBFwZaVfsZGTOn5zN8MeU5rGern/kAVRETQam/YTOF7GG
O0ijDkWqkKQByGBsy9rHv/+dsKO1C0LV9eGBtjh3Xd7rWbImTOAVtK2f5HEj2RserzfrnKD7AB42
xpOrpvcy3oJ5X6zpyVlIbYMQD/NU5Re288sEsNifVToyig8zkoDhxrU6UUc65j1sszaryLeF4Adt
UscqRq2soqHcJRjZzJa+L+TdcnQG9AUt28NIsKbfeyvFMjmKLZs8c1JybyjWwjsKX1RyV5OlMxQI
U1cQf9xvs5RSzGWaAYtgl+q/GL8Rdj0CfGmwCsn4yGiGBQEdkxH4DIYQUbLXgjpDGFX+BbbQslf+
rMEiQsJIi+VpEX254NRXOYge+mrv6tbdCYz9EZjOmbWTgJs6LuqmqNJmOr5Eqt5ptn8OHkk2i1lK
wt+GejeXzqtjR+nfTbFhHqDBwpPgCevpQ2QoWTl+gpRuy520gEgYl4nAslBmm4pbNaPVmiSVGArr
dGt892hisMgDpJM8xvaXFLoaq5BEAet4/6XXwGXVTi+YktAP70CzSZVZYOjFZDODrImMTXsYKim2
YBQSPjsxI2riGc80iZ5uEMIQHQCO6uWNEnVRiq7qvNVUxJmTL9mQj/l2ExDwLAh6t+YZPPt9xhYy
OcBK/Esr7UZBWxNbgsaukVXjssm5Ry9ALUPfrqbssSqyB1zCHYH0lLmDkO3NIyruuFvE9QYy/t/o
EPkkByLXGZAqhIt4DN0imKU40HmDrCyeuzg1YCIeygc7c6gnC2jwrqyJzN4kIxtrMBvUjWEPowms
atN+jIAxBiozn/aKIjl+X2U2Rp8T3GvGdm8/O/Bz842V683KICn+IVeCWyCOjpowbdQZ1LGIYsOq
JXTYWad0sY5LnoQ/DPsMLdqCBaRPO5rIflLhN+WzEWEsXFR9FjbO9O48Iv/FF7fDeVngJ7O1dUvW
QOlp1grqHbpcKmikda+WPR1T8QbLWVq17mDd85zDJmhc4rga+U7JcLekR66EGI68VG3b18EOpuqP
SaYBGrio6ifjxstVhJSav7OL67qJR1BTFCG9PDT0IlIrs2lQTNmzhNZOb+FRysHgE27UkJnn9V9C
FfqJFaLzwRqnH5EZBPslZwykLNqBqEkZjRDEGOfj8fgEAVaDHZ39oL5eRepn43Ub1IT7D+TLfzbc
tNuzxCzz0LjnHG0PMdVUFDccfQnEWyEJmRYs0LOrw+9Gvrf7z4FPxH960IPhWjgG8ddejdTIDZxg
L9lF1djrXpr5cdh+2O9D7Lk6HWxLmXDQ7y0OqVaz2IMH7iDh3ceWq6pXjk72DGZG/5tWNkemTgYu
Ja3iKf6bCpBJbI4WJeTcEI/xO9vmvpSnoHIm+H0la3KQhqdds0vxLCBmSjQ45zyMhedquWAvlL6F
Tofw7tC6Drgz9z88ag0xzsEnKNc1qa3IEod4P/uQ0BlkT8H939IEDT1nDIf1w9F2WINHFQ+icKmk
3od5GwmiBAgkoMpoyoHUtM1IDx+HYY1W9nd8lYWLgb9aqFTZuSCpltbfEsPs80UTPG2yO9M/OP9N
v4dHe7W9dJPRHsI9N6u8jdk6lLiJcY8PeXhwwZ69qhnkLa3oZne2UEkPE1eFMdrQ13wfVYAbhTNA
7aZdQcUW1VyS7xTROXGYrdWP7xlBsuGVYlbns06PIBYhl8cA842Obsn6KDcy3buahowcRmFFae5O
tyBnl/FBim4u3saYmWXHzLeXXh0RNrbHi20WljBBK1tooxK6bot85GX5mmSQN9gDajyfT5IycL33
MKZ2nqWTf34/OCFHLbHj8+iPix3CyNDFXYtF4HNhAdDtOHofVRdDJLiPWX1VTeoc6OMiAYlfDgAX
/6FbiIdVsc+Acip/DcSzbYOlGpjgZfER3vxw0su2qIwO68aRgtP+r6oJ4HPp9xxRbnTrzBRAx+jx
j3KnfFW9b1kZb0S8u6HsWf/+/dy8eMkdA0t/43v/6f0KBOv6mm1lrKFx81RXYLKSoxboery+q1Ms
PqO8eR5jgykMf/jwTXJRevAio/laHsGOE4a5TiXJtRyuXifyZ/VXmusYH/dLXzI8d3DdPlAX2JlW
gE99EiMvI8NWpt5iLGwzOAnWDEnTsDJgdTHJA/+dlRBvTRdWX71h1xApL0/XYYZGx/pFPhg8yqLR
KyoV94ddYPf3To/gnADi0OY2uRz36tMiUElDLfe6B9IAALo8Bl4+k+W/5IqKiOcPFIguEgCQr3du
7GLDMDh8KRe72mYOZerrN/FQijVRGyxMAZgkVMTe2x8fLMFk8Qq7mXetoQR/+u7c5NTflzsDdH9Y
9LtcdOhHAQ8+5B/tT0Q8LEC/B+eNLpFfcznRsw13jrLwknNjBEUP+8mFjaP7uvUNX/JzpMgDHQ/e
UJ8EY82RJHNpmSXvhvG+fCCMWgKlAi5l6vtzMZJ8ZQciwTaj7TXu0l4kkG/ukaUtLu98zIc+0Aa4
/wiCWI26fs8tXKKI2VChZdgOU9gTWYd/+BlgxLq9O3+hw5djFbZRGjfvDtNQqPlBGCej4jafKJuN
vKodY197e//BUcXyCksPZGRW05PWicnWm4urcPcUYBGPgKdkN4x1sR4zQX5zAOBNdWdrb3/NBFLK
MNdUXVfz20puoxDNZGe2OSHPEAY4j93/QbV7Hjrj/caCYIFP4u06QzIYnXbr9l94ZJrEI/QMjKfo
nZf4FgIHikeAkNKBmBUiIeeJFf7gT87SoaRrVuHWx662WMMEA0E9UpeHRMh8gCFbYWXXd1Bj1J2Y
nwx0Vy4jL741cD31BHxJtKsITx5fpbxpD2KReCVS41HgGaKv+JXAuc7wEZIWxWXB7dV6YYqzNKCr
6/+GVvdKma8ZomnEzuOasGg+uYOg5m03KMo26uZDzqds2NtYgCjnXnyaFhUMIN1a/uWdNKox3MjO
xix4GiF6VcfC3Y0BcVJtYBB/6A5c3e4EuR0aBXfrlNiv9gq8n7KPoDzT711bj0Lp2fOwduDCQweN
n6K2CRrg0qgaYxOC15dO7wwM52Fg7c/f/M808ViE4PAoXdKAkno9lX+WkIbfIoHjEC9lyXAjj1ND
gw5F3aw4FJYl8x1jq7Ho226IPD20DNU1s+Uf95nmMUMbtrL1oNppM/vbr8LBE2ssvxNLMMCm46mv
/w5naLGBmWh9b45EBY1zX5p8tNWCXoO03nQh0TLtDxGJcNypfoK6MHgtyfW3ybVcZbI/+Y4yolWJ
3FR+pxx3ZDCxILt/+tn9y8SNAtWOhDIDZiL0MFCNPmvyqDHDOiooxQwrgc2VV5E7XPGYZYZ5pLXo
G/I0kjX5+FVwTBv3pC2HrdU9Nc41K1EgEtxyL9P+ehl8twK7cMOKJoh9Z+QGC4hBQ5k6ErWWNgC2
MOoQHdFytTbz3TUQrsZ7W+Tcb4MpdjPJknVa266+XJDwak9tmnPvXSedJsomx5xEixG4uRIy3AQu
b9O1Z75BleMyjsa49JUerL0dtcKlF5aycWuvu4pUW6JjrpV9giT5E0P8l4MQWTxuQL9LaDVMIFic
A4/JFYb6yhqV6J6i7H+n0DU216ACfpxs+RSlaQcv+HEca7exsap/E0ubTKqhoV9OBdzamot75X+j
SPGsMufq6LAkECQMIiJ+ydT1NvYC38xIIX0ObwYbDJbt9cbIoiCL4Il9XJNQZOOQIlwXYEYkddkV
fWClHgDtlQCBF/RCudxF3bb/4MNIDDwUJFl6pfkOPrP1WM0ujfQuZ9/X+sXEqfUvO0WzFfl3WD42
S0BrdAjgJEA7OGtma8oqFxamLEsaNh8+ag4k2HjWQWwyfrTlyT0VdnvqH6EGurbw6FYxhCWTWqtb
LAlFxCwLBWlp7QmKwJYTbu4OqlMocRu7v/C6t5Zvzg0Ba5nZaRYxCMVeNHhb+/JqAeGTMLKdxgt9
DZ8ZQ2QGGkRFqnev5IWBCFS+zhWHKtLFZW8jHvSQfgRzedhoWixNH2KuZFtmDIhCoFrlxXgUm9bf
QuA8Eef/zYNdXv1LU5fQaxRdZM7mqXEq4oue9+g+nxHxPgOu2Z4t7PxBjhU80T0VNkDB/S0i+E1c
b2uRi5Sp0LokCeg0Tt4yxJRXIWW5N97xweL83w2RErlgamlvn/HUmbSL8n9wW4tf1FL/DDMXqpBo
F3LumK9G33gap/xW1r62M5T/GpiuCT6+sBJJPlZVNckfrFhn7VI7kUDXBEynLhW5dGpDxDJ31nZQ
LD2+K8xpTURaT7pxHwCXOrFEpC8bNt9bb1cooyO//UVJRRcUXYijuKD5Ju3tRaaOt9gf7IspmPyj
nj+YeEb+ZmtEKRLszKxMvd7abBnstN9g9CVlMo6b2khBYg/c6le9OoixKT0emNqSK/JDlOlbBlHX
AbdtPj0urwkFcflKIRzLAEFnj5VPSeN13fmNlZySbyW8doas7/lT9N3dRxub/09qUaTBlhGVLLR/
SyZA/8coC7+uFAdDsDSsjothtPLERiakqQq8Et3qPNB6pZR57z64VimqBaWtfSsQEN5yWWoG6VXG
o/FylvJI5W+adksDRxKEuxn+Xx53y4rzfmran004D2rl8Wkyy4cDi+ROkD2/SLKGT3v8cpnsWID7
PAvxHImI8BtblIyiR1LSpkYIe0srKu1m4Je4bnoTNmpN8ces2KcC9v6d9YBQ5CxbfYMU2Ttj3FS4
cB5T/5YHL5aGTv45jrY7Maz+9fIQ17Vozij4tS9PlXq9fUQFfl6tzMl79nfMIQh2Vev08nYxeT7R
lnWdGHYhmisaW0DCpnzdPILHoCzC5sBwKot+X1ajfN74jB2Zj4I02all3nt+zSwioGUiG9ZvhL9H
D+SO3hQIUAsj/lRUnZT2Nuyqggfc4pAmhhpx/dMw7BI33/Y1G0K6jmMRtNx3tcOPVuN0YNrqgkH3
Hbfq8AsmwqTRI5DWIqIC1vJ0HN/PR26X2yuDO5JDSM84I2iEl1DuXPsJJhLcuyV/yJOgp/GBlocw
2iNNvph1dmsXLDZJORE4UZftzeGwlPeM9cHrjxaS45ymTnGkxPE99+MR5OnrUgbbNsZHnZ6/58KH
1cGOkvZKoWWTUDrdYwwpBjW8XMCD/8pJXudDkQxyA2rC3Rg2A6KJIM0/udPrHD6NDfiH4Aa+HuZ9
6jufnFqerwADY1KJbv2yjV+/ZGKm/6E8JGreM+OE9bVw+8I768FqRwZSi9JQLFuNHvBZwU8tCxMQ
Hh+FXflK/vp34+1zbSqy8Osg5Nw9BY34uSQa+jMonl36iHkCxVEF8B0uBegfOUuItUAoAtgIv1xy
LqiDPuWal1DHVP+7kJr1C5/5nI5tGsZBAOYifKHgEFpf/GdtaB10kwjCowGOfgDa6fkiIvqSaAW5
Y2qdlBLmLOGJOCHODKo60Yr7Kho0xlzAhfAKWfjImOShbAi+U0JIrbEq9I0FDjMEVWYzB7dIT0YZ
29AH8oNAH+Px2Q6q8av9kbr4ftr9Um6QqFJcCqvBXNesimEdoSuoIp0aNtBNqnTA4E3TBockpiSx
gQq2B9ZGg9mOAIL4wivKVYE+zoypPIK4R1H5WBr7Ceh6VbX3glzxXz6qC4F02xjia6G1cMqZFNXQ
mqHqG3AxBcrJIAW3KaAOLw+FiPACNmOz/HVFq8UauKonSEdF7KytG3xY96cAosJfCP1UGeISk1bJ
wxEtwTg7mB8trEesZKPl9kB0PwDQiaCHmF4ZvmSe8DtbEdC3CjbDzq/i1bMUjmJHP11zRZm6Wmsi
h6DWGFCIg4yxrNlt3OXAm3/hF8ENOzlRwIA1MEUvDMnl16ZkkTuJF4iW9/o0B+IYx6Qt9bduj+H6
ZLRzBLMXhZcfqIsI4T00pPkqgCXOI12IPeVKnsV6E+F4g9+qqrXTZ9AWFolCYGLo4v+cmk3G3ExR
et3iFGQci+BakKc6ho/q5YNqf+sbE14iTZGgPzrkNWQ5ea3kuA1agmZ7n94KAHl2i0Z7xJdpcQW2
dx1/iz06Nuvqtb5G4lmPvFVAlghNdXsJCWcPVgJWvodgIH1VMJm/fVvqJSf0zcqgNH59FW7HqI+P
asuZjEvG5cO9blq++4UVAUo3X/710ZrDf7z9syK84uNggCoVW2TfNz40dUN4KIYQPIJAUdami7fc
+m/MaNmsO2Q4bS/h1ULye11uWIuYbKnx54/+QLC0FxD7Kbau/zeKFouZ3oGZywdDws4Hh8pu+wdA
ccOg7LnY8+xaorZa6XRIBz643PkfREsNrEGbPbo576LbakNy0RYeVoCjbhYJ8JfI7O3J/zRSASKG
o+fmAS4PMgcdccMSPlps7fNjhZnJBdxolb0LuzpkUedetFzVMsWDsF6QxCM2SgSwmBlm5h2ASfRH
OCogdVyGMSJOPcW6AnFRcAdvTDk4gDygsN+YQiL+8W5Hd/arn1Y4ZmmlqSJGGp/GasufS8VQS6qV
yqKrbEEUOG+41rGJyQPer/YlAJs15PX4dQmFkVsq2PtZUgk7nUm2qoAlh/AWZKviz8L0pNXvJkgD
vjuz5BuX1dk6LD8MhIIvDJBFWmJH3Dzwd5Ejq21IOFuJYfHpL80VVLPYoLPIHGxi0GdlU0j5f6rt
F3pXW1gey2M/s2T6imsoDokF9s5dk5PchgB+9alVNsHUrRg9lq0dlkPnithB2NAd093bgS6Wo0wX
3BKoO8B4v1NJV0WymxqyZhx1yWTvidZrEKbY9ihpP8MA39de6Zp3Ya8yQCpYidxSqa8phTXIQyX3
w1+nW9cnYdZ1hlUpZfFMDD0+SolJnTjjv5OgCotPePnwMED7099zo3W2FgubaxDTUU00R5Okmakj
GQ1GKXN00nDfDGRmA83q7E5F1iNwRiweQ6om4KojoJWehaIIi0pwAIDKLfbb6Xkc6qamphGcCyI+
FK6BseuoUMF1Kz9orgPVgMMoyhRaNSSaecav1eKpB+AMxnue5WW7VJAsx2VWcC89lWio3bAdmKah
R9uKTjiHtmUxAacQmfqJShXbiLu3a5lUdkXjt3FrLLa1ot6guVID1YNWYZK5MyVswoxWRTUpk+Fr
7/jy0GCyU9XsW+xhKiCerB7tBT8DMN/5sHo12TajHOUphyX3z7WyQ01n7AxabA5Cm7aWFSBQ4itK
nvF7bj//BCMDeOsrdCwPcHJUK0h/jAi+Uv52aF5nedEImSMD9KfuwD6lXdw3KdrWflB3BhvkZIol
pOP1ieAG19AtlLjY6Na31mWW01DaH3gZXY9WWWBHGFkl6i4jrhllz5+sVi0RaMWTUpgwmi01DsHw
XjrrLnIj3tRGckc1SlRspDTsXD0QFhM8YH8h5usTnKbCLmG2h/9/dbncsXkZY4dDfN0uIGTvRGih
bQhcvkrQpJRrS7zmC1wyUlLj7cMKjvoLeYqjJrZGC7hDfuoFxLOMprwjRHPj0YjpgA9M7jyhHhll
A1kHXWI19pOYwd4cCiRbty6HUGjLzADkMocFUONcPI1rIfQK539A12iZc6nYy0G6/3h05OIp4/GW
7rShcM9HlwIiFieB2KCoRa7SqhxVdWdsD95tNY0ikBOg8JMibu1mWTwL08gqu2jox7J6XBTcd+oo
eikvNt0Lb6DOMUbYD0xcSYiINSqHsvo1xb0xPlLJkhxpTOLUrD5oQIBYQsfJFWGtN2saIuVpK0Uk
3pnbHpuKT1oStKwWgw3phn+8XkZiDVtSlkLS6rd81EGpVj2w8tVqAYFw7eWN0pmXKczbr6zSE1CT
rZJIDsL7JXLHGy+N7Q+em52f/6uf2mn8z8o5JpMBiEnvaWOfh5RVqqEWd5h1VmwEJL3ExnrR8ctY
4Em/2XqZlKkqFJmYztHR5Pq9q43LViGRNRPk/ADKCB/G0Nr/TMkchRVBiHiSBkhL9aU0ZmJXmby9
da+Juqlshnnx1ukrO23DznuSMRqiCX6Ncj1tEth812kOu/rtGB1QAAM2FnpW3Rx/+FFQ4EhpekR7
xiQaHzFEkGwRldA4A8zyzVZOdELm+4GZroTrvIteQefu5JE0aDZa1svuC+I2PTvMP79OqdgeeafY
lIcj+Q4dxjng7kpLbvrGU2ETr87tWPA8l8kU+3X0xAps89DD1d0SHQtJV3X3d51iSRGefPf71ZLP
rvnCkZtEZ7OmLwfxLkOgJkZ53G60Xb7Y3HZtR2X7EWkf1tquURH7CduJF2CQjVUlv2oOYcU9Dk6b
AWgVPpfZJWe5pG6aXTDTvjqWTR+xkTTkSDc1AvXw1r1leWI/RkA2Zgef96+eXS6vTTj9cEGJ+IHw
Znz98GYgTMYA5Esym4yRaq20p43DT2VTGkgNV6Kku/csVD1fqwnDqsbtsCoZeATdmdFDSM1Zhm+h
FexcwhaRP4dkL4MDyEbZlEIEeP+rgnHo0M4/514zIwMlW/ddDiCznx1StJ8dUhdT1yfIf7nsmx27
0bvXLcb0qKi3A5+JRcRjtjQdwPHS7/bGpUJ02ytSKxDHw4eVh0/up4UME87RlIdDV1KGO2noY/Oc
zOPEh+/S1jp6OBfhKlAZXwT5SdTpcTmuJo2GoGtx2rlzRgkuPheB/KL+GDhYkE0Tx77XS5cMaAO/
TGHjV3bOa2REK7Ey0wVott94HW3dzXrhuDqk7GFBc9+YlfSdYd2I8iZC+Qd5CwDULkxoO2XW/CkO
kJArZBmtELk2RKKYTEMDUDjJSY0dr5u/rOqoonCGynzI1mFwNT8UC2hfqFD9xw1ZquhqpaxXwQ/w
TBKIaiNnXegJyC768rMx+42chDwico8j6cHOciwc8+qWMnd4Pt7xdASBSMHxPGsLX2K+VUx6Zlue
q8O/HkPyyX0lDFTbPNz3lejCAeAIrtl8gn3L+hONfsTMlNbZPHMboc7t8CIpsE90nxgnXNvGvbEb
Uxa6y5IrOIValiH4a9dTXhteyI9zoYDwjm2S2NnAhm/H+/3Npni7WpW5bMvkg1WCzZ/2BQW3oOqv
a5oZ9iJw2EaPmPIzPiwu7QTT4cVcv4efu6BTzqjSNLpYci1f9xgno9GXxEE6+16rqFUC9TlJ9bqi
dc6cM595Q6WPMDgOM/qwWNUag7L5m8GH1/IkwHeNHpcC49QzSsnC35FjRnFlv3dof4LtboYsJZsA
BHnykjMILhSktZDe2r7v6zsOKnMlg6Svx/9v0UHMQHWrq9r6tj/sCCg8pmckNr/MXUWnE2cegwer
ICn4E2xB6GCbYSNAre7AGkdxvhBr30PvcgqowtANQ88xpGoqnTfknaP2ai8i46QJpsubkvDmK7bY
HamAGX7HS8lNbFtg/Suo3sjxCD7T7zgjpRQpZpyjHUK6oemsviejMtpaOMCelG5Om3RNS2gLh08u
XUqBaIUmvp4iFQNDX3Zj8hExuP2PGtAaPTxReme4hOspa0OBkLjkxTCgEmjs10TRdQSRx1QLqMMx
9hLpOUpIUkmP/MSqY/kJVirXOIGTRJEKIowWraC6dBmLJUwNTBBMCBD1C42WjpOqYWoG0uRbQfZa
SosYRnYGUdOYZTA0zJpqNn4C3AsDBu4x41ePhU4timSyDXUOMis1KK1vgM3VJdKg3U629+wFCDRX
sY5V/FEkA1MmX4b11Woo/wq2boq+t3U3r6HWhYom644NQQDBC+s73eFdvkKPFWKE3lv5ihXZgRgI
cRWjwUb08L7BdfH6iwC8r0Z60JroDJpLH2ri5F6PM0HVC+5o66yHX1LOk3Ckm7mC8Mc+AovXEVIm
LfAN0outBByo7z4tqLiyFGKQQZSzDRoQjm4NINuRwVKtNdZ++FRQmk4T1ksiCzHgF8JDfkBOYtPN
0H6dJQmQkhpmEobm9Pwz5Npsja3CTeoYPBsdHTUftF7ZRLGtzuOSGXl/7SpaNGLJLevCqCzXNBP8
ZVmUOK4G4loa1J39TLuqbPcwjXamMyymWS913gQDOPnqjPP5ipzWIZ7TqZTnk0K8tV1cnJi6xxTr
dXiknbO81/TrCMeu+ZVr6E0B4kFYjuKwGLW5fgY94FPzUiP/svLOIcXn8QwfCMf9y8UXS1gS02++
WJfKDKFl8zyop/62DT3RS4gpEkBreT24U1Cz0XvTXln/V1cvKGpQHbCEPSOpnS+w3QBkWbdQYrjM
jFdsIH1kxFZ3wSzWeS2mzlNkFm1h4cdNeydgkGw0vW4ZInds6Ltscn6wlcyo0PBDqMqeuBf+NuHp
8v/ahP2hYtwTCkHu0PmDAa+8FEgsR0WBGJ/uVxfx/qDzKRbSlS061szLx8F0lQVMnTD5yS/sjXqt
emrCKXX+cVTbvR/o0vQX2Qt7hl61ajtMesEwPDSbolfSNmDTsjG+MVt40IclbPyUErQJv7jVm+E0
L8dJIoM/ABiCwj2a2vdioyr4T6sa0Y5ZKH3foGHcYASloGaFk+iZ92GDopE+8ZmXA2FrayOsEtdW
JXnan9WSM9EKj6xyyGQKREglesZT0NDgQG/bzE5ic4uH4jrw7wSumjQQOFkmFakzj0MkiiPCaX9G
d+blp0DjZpRB8j1tXeSCgw1MW263HudkUnUg9X5QbSlFmR40/j3sLDbm3arWI1T+1Hck/vIjNE3S
88fNjyby+9cojJ4dRB+SYDEocRmdz6j/0IKBUmAQEylEyV2JPWc20KZrcBScE/4w/nZVrOVfYHiG
xGbo93yhsWA9t6VPJ8k8DKECdEBwVe+5f3Ui4CePEyOshSBfxb8Ojg7c630ueiDwjWlGrNhnVqSY
PqR/yjfJvfNiKeKfl34o8FNwH4YzPb/YCpQVph4gyKq9+e9FJ8yETX1TPMokQFeyexG4g8eGvRkP
tKSuT2zaoKiRleCcjX2ZpdQFS0VPHfcXHfduom5ztAC8Wg6f8Z6qwJ8PR+beN7ma0CA5wP5Qy3sJ
cOsnupW14hr2GJKswXJ4JTbr5KIWC7dEXFhhT6iz0UaF7ojLkfPzQ4jLrimXVzdU2iId5CFrkBn3
ZV1TYOnK7niPaNxYZzIeXL4aV2CZF6WatD3/Nrt6DlImhrhyl38DsdXFNSWZjrnGa4HIHBv2+GZm
g3DoTlUEBIgJ6sDI8WYmGAiPUe7u+5YWkbOg+0LiXdnnrubDl4o0k9+h6kat0n8OOh+FuOy3an7p
2T8WKsnkSZvg24vchTV00+k42Cy/HJUISPLjmOTTy9AXquGCCBDDcOdwuwotx1yLQPEWdF//xdBt
/4+8kidMsLZ1YPqSWAZJfA1prGMunE9ZBXUmHkWWT825WfX2sxZby8PL9SfBXs0LbxZZM4tadsXE
jX7bN4fE48khRuLM8SOvsaM6AvzGY15Zakzjo/WDHXbaWI70pAr+8La/8qOgIomJ85hx2Baroxqv
2SdkIQFW5Q6SC8m9VxU8DyPs74QAQQZHqY6GnyI41lBg6xVqgpgnC8SF0tbAGAHRzWvbA6Dxy0qL
nUFq3ZKzlq04MzK1BJIMDLG6ViR8+F6MoQYEuZ+xiPW++oOtpvIp4vBwbvCvKNqADq1q1woQ7ZG8
vwH9trNkG0gYQHe6YMqil9rSxdO5J9XfUZ+yVuJAzbWrzBp6A2drt5Uaj7BLFs5+/Lpw8bFbHNws
couQ9ZT6bLmXIKJbPXUmOWyCRxp0VcBC5ZUHZQXOTFf9qivRSPzB2PRWfIOXM3tyak608kOAb+7b
JOyTNlenC7ZAbVGA8d0Lg8/Q2e29GFClCjgMW6TlPcTQCulz9XWc8mHaA+QzA6BLYFYcG+uUDf/b
WyzmXTyPRl17WfWbHkZkTFLxnCyNpzAVB/6BSR+7TDZWK7cvVZ9fMB7kpjw7OhzrAbPGC1+7wrCM
DjO2or6ptJJcUFpF/g5bONauT/nqnQj6IjFHMwR9XtLZeT9Y0P43ckGtAy7yMdPGZoytLd0MKUlI
vXwUWY08oSqQ91BJYBDb3mdYFz0QFmJypyRO/ktW6rv0AiASR4SJqLSGEnWOD+AU26xYiCCOG9wQ
MW//6u43YQUUK4B6v0HP3GmVyJdA+VL28g7ZPA0ZqiazXwYQ2Envy/mwV1SRSiGRDjzNDRy+5roF
5Wy4GwSH/pOrxLPHy06lNl020J1rBR1LDJfIHG85c32fe2XPDCfPaqbR/4LcoBMMItKvmagxDNvH
BpOC8V665xytNn+AafNjgIW4GxRuUkPBywgwNVxlJzQAdVedddvmmhRDmkiB/NYZVGMLmeymbmr/
YkfoL156md2Sz06CXpUOF3xatqyVwYlafonddjLeQRgDep0IFis3YplInPCX4l5jTYvuJdqsTuyU
j9F+aXhnp4M1dIhkGrGpcbrNOCbVjwTL3ppq1ZDYC3m0qtrL8quYB3M1yb7dNJvuD0y25zK/1sQI
vIo5roxgSa4Y79b7QBG++HjiTFIeFFLxEFuXbIxWNohhS3EPjp9N/J3HgKH7w2kgGAM57wVYWhag
ihZLgcsBozt7XO6clzWSdL73j3DudSL5HD7MUTrlm8DAw5NVdthb7D4Q7/2+BY0igVXlOA5ku+my
zDMawcP/G3BsnedNgC4B5AH/2s4Rze9ynLPGACGMLIDV9sOg4UYOpW0GKCy9yiCtvOrX3AyTcAjN
VWBRoztI65/kBTt0L8IvvUKMJTf7bTGmYCl7QBYmqnSFLGmvlYAh++u6eB5D/jj0YTLnLSD8r+Nz
a4VN9Y+JE1ZMLou0pfz+GxOIiD7eYPuTQ9AlpuH3hjwPCNMyYr9kQiOyg9j0Qw3Oe1kuNYNUt9/T
UYxKPAvzY1MGBnh3MFwfDDt//ujU1+D3/TuYUN4z/fPG/4sheE/CUxR5gsoQgbh7VcILeWwOzggA
EoFa8xgaq+ZO2iirxjGrgW27gGSUNQdMWG8ivbLS+SFjppcgkog8EXFSOWIYkp8fjrKnJ2kECqKN
07Ri+EMzFxF+PjGmjgCb13kUr/Xt09uqnZwndvv+bYjt32Iso38etU/lJw4y1UTCEL2hf9mikUzl
ifZjzME4vmQJEy24PI9W4hggrLDhUtAnbz6dsKaMJjycpSTm1naOVmK7MzD/NOzEDX0cxPgUluI0
bB4x9vzUe7C882YG9fABQ6/qfiMIDKbDgexQML707YVd/WkaPpg+tJG2Cp/dSuJvoeeC1YY4qvIk
4+e1j8NvykumqCYU3Wk2+rcN1WcnECiQfaTrwS4sUBuspDr29oWzMsWFFH3cAORfhDcGM3fm5eVO
SUbJ7IaiQaMI3L8h7Q/M747awX9fRU+0v6uDIr4dB8lc5kdL32wr1Ux4/MgTMpZ6hGWSzXEBz0E4
jTKCVjyTvkYtfHhAThyf5rw5PI0r5AbOcD/mF4MfPAu4ESZyWwS3xtCVjiyXN/o0VYRqN0hubpTy
iaOk7Vl3jbQO16YXFDJeGxy3yQWFSooiw+ayEkWrza4nFnOBSgsu9wEB4zDjltkywMhmxltzXjVb
0m//fWJOkwMc0RygHsbndlAax3NUt/RjRUQy50KK3AcA2+69J/oI/U0nQPaw3X6T5NqqDVeSDbu2
fuPfcDemDAGa3+SmW7NM74WwyOzB5cqKkuPG/hF/lt1+RH04/wId5L00uSNkwIRXBWy8q0Dg+veH
EnAs+fH3Zjb0tsvjQf+oQb0l5ddzdJS69xKOZ7AOy86Z8T3MWWPI0jwn7CrqXdvUTRMIcpy4bcD+
mWoWbUUs5sp3llxY2vcTZHtU2FJi5hJiplWePl9nBcUHjS8GkZPAwLTOMojGD6X36w1XM6+Z8cx7
lqci/2ty8SFvMInM2sgZvQt4ZxL/1F0Giooa1xtozorjeRqc0ZusDJ2/MKvaIcynMnrJFSK1cwT0
7IYSLFyQU/UtZcshGzCF0jP8ZAE6Ihw6u0L8FRU2NcIdNCAHA9aJNKF2Pz8Hz1pQD0PMlInIEF0d
PFY/lCgLMP6+HGL/ldVxFtj6tL3YZTLLH7j/Za88wqZiT3tIGb6LBgS3fEp5BElba0jZboKns+Wg
0IbFxznOpos/ZtAEY01VS1tJi3X9xbY1+L6PVX5PktjoJP07XzIPvQIigFEwEIonXKno4PpQB6YP
EN7GafiOS1CjSI8ocZsSD1rOK5UlPmIpoDFs6D5XWbbVMbvE7G+00KLJQ0fZzfydDOVQqgOdx2Tw
eltrdoASLgI1eUD1J1Qwet64iHpAfIFTXdNwHOda5XGJXh85k59Rk9C3Sk4Q/FLJwmadms7ehEfL
w6Li5RscTGfDZ6nvhfQ+xiQtT95vugdNKIhOcE+5w5fzouNq/mkME2W3TscaX2zsXv28OEzopMEm
LqX8n1VMzohyOWXr75T6Me5bgl/zYtuqjl420vgyp2ozLv/QPu2VApXLsvuKlBiEXfwnQaZMrDMe
mXOmY1thlsyOTEvm8PdNvGjClOzifgNkTIVVzP2CAufSG/E41rSQsx6LZszCdvIeErmUP3ofkUYt
3guiyfMS2nyp1jTHHhtlCXucjhKZ1EF0ioqlY3HtG/HHxC2qHukptnxHYSgkrnt52K9wRtHfE17s
8nWlCbDrRYSxF7gxDjeTo9xT+UzzsI/CNOLV8jPIi6ui0nkvwp9G9XC5ZOV10euQwc6LUn0Njffi
fOFcNv36HfAwex4roabXbRMwyGsllhTtTq2oOfMHDugveEfmBxWGuq4l1p5z/gyIRHgTXL2KtGfF
M5t5KFkm2+xwnSuxhTD6KQHTz/0zWTFurtvHp08OPzftjXhrqmfnerxPeP5Z/YI3zg0XuY8P6VJ8
4aaA6cJn1OGlYdoBFSxQxRz1YbT1WW1yKYGkLGJ8qBqbdf/x3G1iatwGQxlV53PJbwcE9ZmZ1RXu
h8yLMiGWgnColmH7ZAPNnUgMvYQ5d4jmJVx6EMnQTxF49dIwlQ+QPGY838qMciSmrjhIO/wTfZw1
Cd7NJ4EsDT3u76Ql2v28xEZPlbVN7kJZEWxjZVXrbaSwbs2bK4HVyMy46G0afriYzaCaf8qHHosZ
JKeL1XuuhhPVkUZ/zt8aCSkM8qn14ilON3A2coHPaA+1aaM8MSKgmEk3WwcX/YFbM67e0O8pOT/4
c/Cq09yt799Gbi10eFxBCd4xk7KX4qATe7nljG0cio/zP+0h6VbSKvvVthx4haWZO3DglLjJVaiJ
FzJPhdCn8Fyr/n9NrN4CM/cRR66BcWAQwk9F1SmA1RGLVQZ/eUhee+au5kCxPdv5/5PgCJsnDaYN
Eeq4bIKtwYyJXFZ2BULWk1UxsG0FfDnRnxM6gufbRX3AV4Xaj1FqFciMsU9vFKemF+ymgr34M7cV
uXLZpyfCDjFAoUJ1a0oOrXKZrJ3inDh3nG0vpG6pYlsFnSdTyKd56EuOvhZIIqQfs+kSAqcfu9tv
wR+lQ66qfYtMRgDyms+GVCibOXoVvU5VbF2hnxwZtxNeFVNddBGc1GuoFLAyMoSAHCxULu6zzMQX
AV6WLY4G/CK8R1/3MyopnOx9GKsf0jNldnZA9+Z9v2NHXoUs6+lAwWJ2NWthjFcvPKwM0YL+epuw
hG62xJ7UDgAwQPUOdT6wX8zp+HET7YWYZS+DtPzxrM/NKWE/xo8ZqFMP5WCtjLBouYHiTLp6Nf3d
60m/g4sCbMk9vnoyomK8jIXBmxOEgPB4JsAeaROkt77ZKhWCWgidz2D5GtfwevU6mMB0FVh/3IQT
0ugkBuDmphIBwwAy4y3gZ7fQ/WPKyzaBAPFZMr68sJVMlervXoZRmPUj5WwEKE83p615/ahZ4yfY
Fe8jwwWJFvnTLnxbrSFJlTFOJ3dOp5lsDuOp2djvcI/L7hApst1Yq9ksr1fJ0im/TJ9BHHBJ8aZz
qIycddvM/qth3OgKv4H2aHKq/d0zguxk7+4QXhCG7b4l2HeNzz5VdBUOdBhAP/hpVr2ZadH9jCRA
LTOYGzq4utNAUKARwZFyjGptUFXj4VzvtZB93lSTltpkfES6Ssr7uXkRTRQui7X3cMAq05riIN3i
L1faTRJllSeple45HM8w+sC/E0RAmoDZsnNvunE47yLRc+2evShzzSQAv4d2bOzA3EHOPQuvKvJy
eO8bM9tgJxkeT/er7Gns253S6p+uh9Qy3WgivNcR6yoThKrFlrw7gYmGZ3ztrFTw73MMshPDN+vc
hSBuv2s5AslnSm4+iRMsuBu9mg6C9SH81GbDYWuMmtqDpmdpep6H/s73ohFMFEUjwk7eR5+04JUp
cIu4wsbcM1GilCqITVB9xiHH5nT7qDKgo9qPTOE8JXbwljBhYLkSIead9BlLITnUeswj9uVEcy8y
n/9VatyDGN5GjUeSvua5IDYVpP+/eQ30HsvEqeOH4082HrABvjfMW1J1kuF6m/2Jts3PHHxLY9gy
j9jFmzS7vCUk2+2MTa/4ITeJaGidm4RoRhwhVqKAA7mLgg87ki6bONDDg8HjGO8YSeixmNa2JKmR
DDJmtJWrtqlDodirYx2S0OHK/tTG2IPrzoliT3QLvv6r+rNZqRImWKgiMHCFEs8M63bYriBvBzM9
D9BQVFNwo+JE7bxFBTmEwhia+jsP5fN78472Fopt/Q/7Eakb142D+oc32a8Vvd1SMV/dKAencm3K
QF8IoxYADaQ76icb2GVj2NF8NlMBw7g9g2r1mDG7IQOg8kTYqsM0y06hQ5lhveDL9FkgfumfrhS+
aHv0jVJqmquDbuwGnIByV/7xbTOAGEoGZrkg7ntnKNS8TwMvgHwWJ5rgDtVnxrgWm2sfiBHPAQZ3
gbbd3zFQHeV9SBsvRdFqnGcP9wVY7FDpVoRUYDnr31jvzg5ZwIZFOO6/8LCOCXkTicxID0Yt1ax7
VMh4YV1nclNXBwqcLEPmZ34ZhZJLOLCHeW8tFkDkOgTgO0+1hpDWJs8Y5wzjB5v6+QEPj+JJBQA/
hWHmKwVWYbhknV8D4frA3S6b1SYAOWRm4CgtNp8+MuDVEKFvKAfNEtJS/qTylvguot9bl29VpB6c
XriNebJwsOk1d/2jLMjMvmMq07ML2mn94WolQaf6woi/Rb02YGPkkBocBzA5RvJ6sWuHP5GkouWp
xqm2I/EViCVMt151gT/FuSD1XdNt3WdvityZbtyi0otpog9EYXW35+XJGiqoHmdMOErWvOqKyCYO
4F0s4GFea1blzhqCRcx3/9PeSVnL3xoa7nIN79RlVbcoUebClwmsh6nsbJoFK7tIWFOo/YKgJGIw
xK1FgHxBU0uSghK8k0lMCMka0Kh11N2TXevspBvbvT2ErSbKFovC8HnCKfuRnhn4R9VRZV1JJT+O
M6s6N8+q7FLCN51k8aQ7eFS8MgyXxg9M259xLohqc/Cm7Flwr5FxLLn9v/zE+QBrwxab7Ajt1E4N
9dsgiWvfHVRNT1b3dtYYxR3FiiqzZ+aLinXcKZYxfGfT8XHRIpYRk7NgUNUmVDx6rvwpxOQY5jev
P3PYgnNeZu9IzPZZat0CFoWjW2xQvOXFWQSCRBz9OweCb7gw33KNkOAGTNZBesiIat4JK631i50q
WpYi/1UaWcBh29cuFyAqJuOyk8dEdRktj7RFPaOzOWHvpwPVDaqcOQDGZHft5KxL6LjyoYC/TODQ
1qCIloCzbJh6Ya03dFXSN2E1BomcMKWTx2LM8m6Xja7+Yb/qWmXG/GF6IyRnKxzLnbNtr4f+ydg5
QsL0qn7ns2OKpiRPIkZrydiLdPMsmDaDHHQZrZH3xdO8L+XJ8pGUntvaD+YcMuDZW8xD1Ek8/MpV
G6BdmYVSY/Mj9MwdDcYnXK6IlOqxP0FOG/cSKyl0SJO9Sh6qa79smiRYMAhZVsbdz6EIOJB0Od+x
a09zVsZgnRYfuoljfMZKag1+yM/81IuRBUMIQCqtLFYRyWPMoqYIlWzfzcMjZ+pgdrWNqOriuswS
v7iM8ecXSn2mZT+jFpQWw8IRyzbXVn82dj5FP41aN3wenHUG7nJWtMiHV4SDUJaM9Rk/CQGQbG52
9RlYMG17m64NzI5kxnsOuJX1Oa4pSHDF4zYGXibWGzabu/3mV5F3SyVcn3Wu0wTr5zH6VE34kRwp
dUIhvgydaQYRooC6G7DEVCOs0+gZ0SkOKwNGQncV27OsX9npLw89gG6x5PqdbKNyxOnPfsiyb3Px
1z2IO1GW75TAQ+QBj8BNpnjueNAbKOGnjL1VMHLR4N1+AyTGBoiri3L5P2E8jzx03b3cpOHJrJTQ
n+rJoW2U/g9C9TdZzWJNykpZtRmca1gZtFxQYBGjJpHeF/pHhrtyGDwzWhJ1w+wGyhg47JP2ZV8y
ypV80XePrGxWaG+CoowcITS0iNs4nEOkKzoGixRk6YW5gB3pNpe44Ycdx1vjNav2R93RH2NzK4rJ
TgT3ICJeA+kr/G1MPAMmThjrOARJ29BT87Pq41go/m5tJITtTlbc8z/qHpoKGO8fJUMzOc9MaG55
hlB0H6rvorXdC6mzS2uvV457h6BfiX6ILz8R0v4hl89DmdBCK9J4SACPOrxp2/sWJw9rs3TfVjW3
8lq8eWPWBCKtVCQzJfozyw8cpVHksGp0b4/HLWpQoVTak9rxCl6yTyjRicYGyweTnzNAnGwKeUJR
VA3YAu5EhoDPsOQFtXcGzLm39mlCq7DEUSt0DTTUBmcTL69Qd5Poo3AxfD+Kxz2V+1W6QdNbV8+U
5YuEOuZHp2FNnoeU6/trNiIs7qq7t8loMVvaROCwJMwI+YM3iK4emH0F4vLJzSFFLZbktUN432YJ
a4b8G5sd5XEXyzRpGxEJx37zoNflA7B+NEBjynk0ys25Nor51TYo49OMWqHe4iE/8oXyxb8xNm+m
WNb2EPvl9jW+mVEEm42l8mBeZMG4pr9XJTZI8XFtmvrbzeebCSZnqdwrSzsAqzVRS+drLWfcNMm+
+QdH9an/WuU4E/AhEi+K1HwlFiTO6Hmyhe1ZYxmq3fSn4lAaf9tL+2mzZ0q85nI1joxhfYPi187W
A5hz6QxNOQDx6QStLTg16NifB7Fiw5PfLoQTensM+YRTNW5nQhLkvZt18E6DR3l7tJKdmN6TU7HH
+IkZv9IrNscNXKLHzfPp95LoFMMJFx6IJ/wE3/DzgXr9EpF+KePvdBa+WxjD8VP1xm/0hxk5x1iQ
Hd9F3Hc9vlSD76prkxQnc91sUea11bhgsrDN2sE4GSb3FbacxscMTP47VdYlxamgYZ5hmtzVfi1c
gkIdAbpjAEzLYG3jE7VOfeRxNwetxpJbhaC3oxX9YjA0vpiwKBfIRenCTfO3Ypl/TyBZENO4z/FV
r0m8SSLNxpGqx3S6u3Rnz7UZPKaeHaTLyGsdGjN8AxQjgJT3HEbWMIizjwdqcQOcaD/rX8ds3XZL
pTcma+yFdY/OEiFXhkHdfABDltgzGWuM4Y2jl73rDaMYIb8z431Fj7EO28ziEPz+prEXlwlVEdy6
6H1E9h31OZKZn++lWAXWnepPc1x7m/leT4SyS/TloDr55lRtyFWas1CqmnGnRwE79kDflDqiy7tm
DD2a8N/r3b3t90EcogP3J+iOIOqKfyLBZGbhpVolmVvBRuAfKCwjtHUJpWdU0Ugc8eBARRYnIxET
zQFDJWNrD3stsVzJcuoeLCLay0UWxZZeUUg2Iet5M9Z19veMxesAit/vveGJAIKBPD42FEMMo0FB
xMKT/e4exf0mklj6809RpuY6yjeW2IvxpwIxv7VcQ7iNiwolAX6Byz54Uouc5Vsi9tQ2JpdsI2Il
4lAzBiBKpUoMYgbxufZQ5sEas20cx8MS6sJHa/QkPPBZ7of5wi99NNBD3L8ffkSKapVAXT7Sq/Kk
aLAxpOncGmwonTRvuZWwbqKd4b3J9BHYncfX/NIr1iD4TQF3ipLSOs+JHDzNW47yc3kxEw//W9i9
bf7Iv+hxxPreG+BtXqyec24svRkboYtlOAjpH1jzZkal8oQX0vxKjHzzmjjW9UWTMYLCxSgbB16c
TfIAqeiDTsed4/JXO/7ivGXGXlORyOmeuLYQOJsTC26KmZA6dbcInrGw6xwcF99MDtsdgGx0FIni
J4RQm1DHsmmyMPj9CGQqNZ1BjTIMaAGds4VKkLUNw+oBicktox/0xOxatekt8g7s3QJd3f22kQUp
MUj4LYUL5f1kV+YHqOl3q2RYyM0n7bnWoowQLRRwSggE++mBOPW3m1m0BNzugGhS8v77pSONOOyI
7icEniHWd6e8/LkzjanahoGcbsWKGC4Ow6amHhamLxvumA/kxk56RzBqmCYrt9Z8rMjL1ktgA71w
qWRdHN+xUCTtlaRx8CtTN7/PgsXfFegPHKdhpEGL/6wW1fB9n4ReN9ZC9KF/NTAnv8e9N9NL6JHF
Xtk49zTQqamT+eTfYGim2EAkRomj1PPbgDMOTurnnDdbucFLKcvJ1X0qs8DO8G4C16JCzQekR40V
4kmxpy83xFuyXMnnaq+W7BGd/2xbaldq1WeDi6BJmSm9cz5v33C1b+cP11IIHi1+nWtOTtTTCoVQ
aPfFjkk3uMP1elemtlGPmYpb95tJxA70hV1WF8AX+nokS/wU1WNyC6vRp9I+NOxDP11P+CMQ0nVu
VI/Jyq5Uha3aDA/8niAb+YN8JCsGnSoxPNGHOJoZ3Lgl5mQGs+/Mb/xtuCf1URLZdoYT14K4D0r3
ROPX2029hooXSGD1xtK3ZeNdYv210erJkADmbBU8JjUNkqyAHim8SmELfbd8EjrAdCg4gAF9gLRv
b/Y6qWucDCtseAKt3G2mN1H6M2ncOz4i2aeHl9pDeBFn3UjfRSsUBEPqGyrXRwNjRumpN/4UQCvg
mCTUiz7J74/9bJ5fLzV3HIUr9h07MlTEtMs440lVUUpBObRko44JNW7EBDaxt6RJMgixShQwMjmG
77kv1hvQlQJz9JVF5OidY9Y5nEZIgLbMkThr2IjYZ4KxNgbQMD0P5fgS/fumwnPiHHh00xham4UJ
t2p4AKeFt5kXioL87ac3Ubml8mAls/F7KiTMxjQtrSm75U6NZZ9EVNUac1eTnfy4vkPBBc9dMBzy
crk9CCxC1IcX9wbIQgSdAtjLjHho1UwyXzrE+hTKjPh01nrvs+km7oskjRf7LCew1x8nj03xw7bC
lD/fM9MbSch7NL1uHaC519x4h6Ne8KOgujD2d9aDeVVmWGnHdC5QIfV4zSoKdJ5nYF3hKr4ysWrR
07+dBvrqJQAD4JSpqKHI7uzguoAD/RX/aL0/hY2PXEQvSBMRG2IdqVWj9y7x4M4SULGGkZqNZWpm
31fiuTXMaMQTI4MKohN3VtNB5O5FUJ/fjMxOpIDjMrHdgjlaCZ5BA5MS/jOjbGjKYHfcRxs59/Cn
FiHqjD0Ivn2SAaNrLU0luqTIXXifyL/PJTZ0r7penx1P3H9+xVdOkdg3UZ1W8gao2Zv33YbElgy/
QRhOcMLSqp7TYMJ2vUUbBdzcCx7+tnYUOQjMjD1jT0VzurYjjkn6+dQCV90RPA4nqxSVzVZu4dGn
HOwhmfV5coPQm8KarIIl23bo7BzGzqmW6IBABfaNmgEHhwncmaVCLvPQgjiNECfrkW1M8HEvvQO7
9JbunelNAKNl7dsBbV+4ilKtC+lB0s7Jn9Wj4dOV/OIOjXQdcduZzPY1V6aSJN9SXD2E5eKvq5rM
EvpKaa7WGGMrJnke2HPllBo8hCYk+ygYYaUyWC+WJIOmZ8V0Lw0ZTpP6sx26Drv9XBwTBJT2WSRr
NVlKMe49oCibYtM4KJRpvmCV9Oew6omhg4kXYrzQ+GNq4fAzDuO1HWUl3SD/vfl4mguVRxR6hdn4
9DkgOwkXk6aMUqRvrxaZRKX6MDXP/5v1Cr8tzJ+xjPD5dCiBXo5Jb9qDp3tcnJsGeFejy0koCGUT
zcAmLsR9g9vzMCBDHUnCL7vkL/kpOoaGJmmxowyk4y4Jkgv00A7716utWcgQyotq7p0sFGA+Kb9e
J0NQlPacTvKe1w/AQHem1peQThd50OEr2qSJApxqcgJQiKwuswPR0gtIl2PfSEUQDWoKF/LSZZST
fqsEJMRMkLP/Cydv5I3So+wsc7RAU/fUNLbuRLtat6m1O4S4LNpwOL5yp29kdf8UyxWyL7hSrxTm
/6azVoRF5lfJrXbZo6xpi7i+N7zl4EM/kFXRFVgL1/vTMHig8Y+9qj72B4hbumYUNpZFuyJwyGVo
PfrBdNfe8ygtPA1V5HfkKa2vZu5mA1wwGbPoCd2X5DRLiCX/e2NSqxH5+sxLhf93FAS3JxD8wayW
Q0zTsWLZfc+cHz8O2/8jguWeDfv3enEsmRGssG3Jgqtx558QX6zEwtdEFq8ysKQ15NqHA88D+1H/
GE8gHib5H65ssmiM8Z0WqZ7kSF1ZD6gp0SF6YtxDqEsaItXXgI4rCBFD9eKT0Eq8KwdQLnnXTqVD
wbMLHNhwimOGDBPt8W46hDW29IgKhRLZcKRO/kb//gLjvBbB8hwaZTSIG3ABfgXLWlUIfnlqVJwU
kCYTXgZ3B2dUWW3iOYDPt5L4PNGn0oOVvC3W17BjIc/vlhVSDynY/NM9ULX+cV8JqguRZg9V2aKv
zj4Abp2BzSIYAEOL2KeWXVYwhlQDXwNNCwM4GUzWrDtI/onpMlncCHSZo89leeTxWtQCZsYtalWN
QD2f+72NqagpDRuT8Zo0hS4/xPo7HsFvi8zpm06n1g5sdDEmiF2O1lrc3P+rEHogPDR5mdbOFsDg
C+0NWJ2WDj8DT5v6n6qskyzJaAsCAHU9IB3dWugudECUUFm3DyTpSrY3o2Fex7jlnXkM+IOqdxvA
mwcioET4aiIO+BHG3lG2PLRGDxioIQRNpkkpVkYX4lSy0T8ZsRZr5vex9q83Y0HOuOJn49c7x3J5
YMQZ5hOBS46q/gHav0C1DUR7XmjPxIAHPQ0z7BOi7t7VlnrVSmBNr054tRCFu1t7dz6iwO1xWP7q
JIx4mwptv40eRm4ZfyiKFLT5BhxCwXE3FhnELTw9tBuV8SQ1zDGwpr4aVLypW/MAUp0u8ElWL9u7
7JDVNtz88IVZi9JXkE4ZhEHpUvmUAwmCtvrTryw2j//QYb8tnWQ+rNQzEE0gFnlUFBOTvb0fdXii
guHcZ/93cEeiy9pwUgnZQOoKOhpi5AUMqLS5zpo/u7HTvRUp3qicv2fIXI4lrDPF1WLNLx18UPDP
YLkW2nE1GEAG7FLkpn2agJ9eZjpWo3mGclIUvku1CFKBFCljZfI053GKpWsNIjBFIw3MRJOWHsg1
cNoQO2UYJyP9ZFA6edrAepTaC4iWZwHbGvc+BWfp3B8eueqLI8Mx6XpMyqIDDy0OFvtGanKZfNlI
/pGuEuTZ0Fvw+B9C1ONPf8FZcmsJ8b09pfTUAjqWY4J1ERgxKzocX8+P2kKyfn/kbsSVPtqFZsDi
JLBLSvOU7aKezYfFRhOIqM1P/ou9k93zkhM5lQozkETv2eHaOZWvAm55aL4+xjLAL9cMhYz6ZvZN
UHww4gyRvi+2tXMFd4q6EyU+gocsmq08uqGeVBgMyoBB3Wg04nBmvJFwgEWQFuVIM5Q51eW36rEJ
/VvcssSygs1YT18qGIpUvzSFrCAMzXwNqHBE8irSMWLslw56Fmon4x36gpmJXP+3HovmhuZHiJqE
SIariqHVkm6lTnpXh3Kg2kvO4QI5BorqGZJ7ODnMwfsrT4FWNh2GifdsfksGJiwn9jT7yyW4vqxO
m7BGj0bNOVb5G2u1mt25/0KxQTPI0/ieOiwnO/CknX3neWAypEndz7sAl+269S2blbiB0MvtaJ5n
JJTJh4G0yv/Z2fT3QvecTjr3VGhdHfwO6l6OmKa5HgaFbFAP93YU5/aaopzT3BsBqoWA6WWpuswM
UBstFq5TRDlHngNCLZi4LoodFmrR5nTfO7o1NVti2zvkPZ9Kdd+EDihyHJwfUOx2z2RVcWNV1A3Q
4qv3vGwGFt5CAF9uj+Ky97l4Om8dH0Csy2WF38Bk2QMMBSrSJ8UYeC6AO2M34Bc/nsFbWYj1GV/s
qVtYU1nDaQ45/u86d7JuZXRTzmPVxuqvTJsRbHzYQuPehoB72pkl1Z7sSSJOUWFz6lfBdNqQgkXA
WIyxrft1ZX38ZV1593uiN8bxW2w5lcURHwoXI3P7xk+OVy8TH9PnDRsKCoSkzFPWAy5KqhZWkf9h
F72zeQYqhj20O5l2czzAEVRdzXKSvFDJRJJrULTxG1BCVqYv9B5DAfRko1mWs1DjBwanSIdo//YK
fedsKgdaq0gytradOiWEXuRTbSxxJnfmTbop1KvViTvDPYyQ28tvaRxH725jMU1S5cHDn0yoULLL
K9B5bASSNOwIJvVZyMPvdFnu1CCJLENbGK5H94uJDDniSdtzQrrWzoeZR3XVfBTEV43k5Aks4EPP
XT+EUmQqzIc7FAXSoDDw7LyiCRM+4zrkRA4Obhr/nyTW1mqgxhlw9G/JFVZbXRUGChu1kEXPQUj9
zUrFZGCrBC4Hy+07vfvLJvchOnTvh1+XqEn5KaZNq/gXg7VV3TgL2m790pgrdyOe16mOshOWc0+Y
p3NOpzcph5bpnuy0OlP3aG0TyiuZsOIAUfFxu6Xuds0MU64RORBG6twO+UXMAMBaPdDZwY+bEEx6
dRHRKv/Ajc83124/Sgxw8FdvCjFiGirX5MDcrCrR7mkLyq26DGJOf7mdSUa09NCEUg/M+6ser6hB
qjmXK/QRLk4GBdDjcWl6n9eIkhse2E14UlS0FjBkr4jJJtdpfOmBOM2j9lsKUjn9z1O38VPhOU59
fpUgW7GRTCMqKxauy0WXhX2ZhoxE7rqkf30zOSxUCi3wiUlDtW+t6t8Yz+pEhxFanZNLAenaRhfa
9fJj7Oq4Cfv8Qjeq/R/c/BFOnOn3tAo8jZumGeiaRJc8ti4KR1z4CuMTQX8D8zvwx9KsN5D+byU9
l0+zmGcAdYFfFMZA/YOnpZHSavtSYkE6HVYokQthFm0LqkmGWJXtr2ZHdJJRtPO4gIe0riZqC0Fr
jkopeMylLpM1IbUGzP3cw0uORhnTJkJKGlgHOjB5G/QsgKGWElO9gpbu0NFcMWu4kK+FcTSruGXE
7jmrum7VKFAJh8j5/pHBD5X3wkMyd769EL5atdlvREIq9AvA9R2E81UV4csC6csQfNazTKfcfPmB
mt3SsFMvcVg9a51GHa0nOnv4rwUu7zdzYM8ELPvYpjKf2XVNWYDoUBdmbgTieMqbyEGm26rfqW1O
ZTBDvt5fLvebBc1gB1L/m52Zg4YDE8mGgNRM02CLGretgqe2w3j7V+2jtpJR74P9deePCPOjWeBU
YYn+hpvTNoChdCz1oQzase0AK7BpK+kh+ouGqqqkhRUnkbSnHrIjNQuFbr6+NVWAhBHA//CoGDIl
CL9ItqMndpPRkvK3/+b/RAoBC54pq9vSH14DegDpkz5lKyN5inKjtq2uT5JOt/AtRS8pVXdw67BO
F8q0IuyaZNiFC3aVsRnaN9DdRfFxSQOQ+8d/rnxQg3WyOd7dxGWSYtJjQeGJ90AGh/GSaOpKJJSC
vY8AZqOwtmUjc04yXHz6uvXHK9KveIa4s45rDdmwmpbhrtPtnIYFWFucZ4/z0iCARDwTGX0VqqTw
t3AHzdwq7wWLKwppZLXKx2HChmQwg2HprsmOQoA5Q9Oa+T19LBD70V4cZmAq5mlJQBW3GALd7Sia
Owe3kcPWvANnpJUOYelY+WdftaUuqGKx9emgG+aInhm9zHb7qX7beDsru9rTcS6VaWEQ0Ew2aTKk
KzXVUvKf+LshIbFXbYo1il5XYRGCin4n0+q6pSPr2+9Oq1dROUxdTpm/0K9EVrqC1BgTPtgabI4I
HN6mqBzewkSyTqOGKwO1MlbTSG6it+TJSic0VVVpRGlKPzLBCrQWWs2icrT63tIxeWkTDMUqPfAX
kTlbUs6hjrnr5fS20eYaGDjEKoWlf0iDZP/r4LblnUiFS/yvkfoGBX7q3QydDRmcwCQLb9oU4bO8
9bGRYyJLaehja9IknchykV+/uCMCowOy+2FE4AW576DxB3+Ubw/ptAHAp4whdMbO8P21u/fXcci9
Mr/FESIgD8nVZtZmG7+hWNtVOFzQp8EDyoU1IXgGJigbRLOAGN5iIa1dY+fDZwJ5e0i2kvwik09x
pRPXrf3jYC6pb2v51gBlYfwE36BMAvTbGyT8Bj1kVdBHp2dTZUE+fPa8ve3M5b4cGYsr16RU4qbj
+mmsnVwsHuUbSgxhUMPSrusYXzfE9LkfXwzGVQAZxqnRwB8fgmS74yQsEXQTlok96yWRNI8N0Nt4
MebvrlXwuN5jBtWTGHdl9oIzEPoOOt3ckPkSoLHfb0cR9WqJKg97q8M2uz0PfZB/2DTQ14oaTEix
j1WAhb09VJIxmd/KnCl2raI7KZ45M8fDJvwCXoNPwQZ6YndN9hyJyncYkhw5RHhTAnAWL18lUJ6+
ET7bvN84L0+/BGrpWpnnQZS0ZZ2Fh32PjVt0WGqfcntpkFkqDhTi5BFSu/GuNVaom884Z8fTU3Y+
6GwFJcfRpvi/pKPMhPeAGsuKz1lC003Tm3EhrCxE/Vgma+13ht9ULEQ4EttE83zYvIBY7aBJ9f9c
h5iLKkeR1kXuIY+L3cB+UVd6jL1o/se/9ZSI9NSPPO0v/acshDt7xFX4UDKCHWJNmRxW8NvRkIbN
SI2RS+OULGoVwdUT5Y8sz5Hsyh6lbDYakmhL4jpwOucmmxAkneF/SlZQuUIxASXciKu5A31BG+Fa
sGQb0/JqSIw5fMTKKpAsnPRwdulEGNotyIF+CFAvPM1DD1BPhTXUgHo9gNlL+JWC0dzh2xQVdOim
OCa4sPTTZe40g04cp7kSMEt7Di8NFkWBTMvpH/JeXJJzoVuLhy2TX3pN1u+p354W9cgCauAkg212
9nowmsB/HFHzR5B+BpXkl4Q3zJwVgUh/56/ZOVECt7dTNv/kRVIzASHEBPcjshsFhIojMK7lDDDr
ddWxOfkYz9fpwWc0SbQOIKF8onpd1BV0BNUMdgQdVmoeenYT7dKdPwHNXJ0Fqpi1Nrc0qeazDDig
WM5eo32GKIaoyH59VUKlI2npSvJwWA2/cCn94TQVfhINjaElxD9pEsyBEBSuNYNwnh6uSK6lwGzV
oM/q8b7odbFEyNWiUisdH8TFH1TgoWsVO2SEfFdh9WiSZOdTzHOjUs1WBdo0Pmg5DEqG7yVdBB41
fdsT+agFBrRJMhkzPaCF7kkfD3/DPgUlXGATXpJMulBd872QXBkkXpGCiuK7QfHnv7IHqGcqzx0g
sj4FCICvech8vRLalb2QIZOXV0IeXMzGStNevG88okbqDsc6db8ve/Gr47BQyX6vdl9275GqoKQk
vWvQFAjwTgPHwy0659SpJO4vxTO82EA/yXKUCORk1PfwCPNNGkQJsFp9Bx+JeOGYMluXREz0Rmmz
I3+h1luMbOgTcupBgPV0qb2r+9F97d22CI8rnrH/u68COfyoemRdbsucR9LlprnBxvM/zVMC8WSa
vnQGfMGCGYTP3FNksDCbzEa6ENFc8vGZIDzX/bz6BamzbWUwTllJ/g8B/6tubNHnUwk3EXDlw2RR
m7quQLoBN8YrF1eSHAA5xYfIz/yhqPinM9tioHrwNb9sus8J58Hz7Oo+HwIol4vx2fRyuyjnYml3
w+Xemjjh3I+QOIaf5uwkYpP49QFzytFBKqAIjwX8seya8WpQkbqPgMgJLmH8uC8iymyge4jNoQzi
fKjIiI+dPVBgFmjz9n+pNJ1Y3QlRe4TuU6d9irq4NI0prnDRBfWbH1xHiGvWr0liftfd5caXAivG
ueF+qsgS9s6RARz95t/mkLtuNNe0rCWeWaiDbeqVWcbJp7DU8yLLOwi/rB4tCm0NLCzbt92wPRhN
u6NMHUftBbTVUOXqf94zskir7G2NWyB8hdj/Sp0N457o2nifiMIY21PB8A4zRS12CHfbAkGYzTn7
hj6vNUGVFGQoeToLYp/nqGB0pZegcYl/7p+QuTxbrbDPo3uTFv1cApTnSXPnQ6Udjn2G+cgCm2+G
piiLV1IxQTPZiZEapsce6iZshJsEnjAL7LejStkeZUcP8BBjb4Z7O54ZXEIZwV4x5now1Rf0PyuF
RQgvEf3j1e9rQzJrB/9lUNoIij0OXuXGDVzAHwuFK9jNMNooun2BbxLiaFIPR5QC+pCQ3NiGp7Qc
slnOKQaLajsD/b7LQ1xstjQ7SEbW13XEfe4VH7tuRdhkFU/tQjEQb0pS5NessDwcJomGXnmxDhe8
EWpDvTNSua42Z7UWY36niPpfQd48twGAlg+hgqeCn3ztqiaCugYhKnA0lAjhSjPZ20Wp9MDZONBY
j6gQGFl2G9gRaubVUJC91iLj9wk+Bqj5Pnac6qDIQmWHGx+sndRAt/wjQn/Me8+NHZS/kj3toVVw
tpP34tOPABHl27nf2TKTx/WDQefqPzIJi50pPyOlK9zAnM7aahX/YNZwCAmNRFPueNx25kCD40Jw
DQQfeBYVNB2DSa7d6vQwahx4iXRoV8x+Cyj1ixrkcZjFxKrmcfoV6Rn19H51VfjWeQiPnfdm6Rgf
CPC7roS0VWP2cbaMlzTTTnG+VIezOpPZKvSgci2lttVTv679xbyJ55df3PULKJU+jdBNuTf9Qcsc
OTMkMmKO+xXv7W+E+nJm+VCcfKL7V8nFOf/5gURITBiOaFFpN43wPtkQbyyXU+aUSwJfTgyj46Yc
2L4VbuMi5ngpAJwib3EnGwjwm3v+g01O0N2If2rYXM4Mkj8Qv3GB/WmQrS5GYwRMsAgfTizoLEAy
xgo96Nfats9zxRNJJ5FMqpEXiNpIkgorti8sFEAeTNrrYihOe6gfHLYq9GgQox6U+UqSz9vkagUl
d2U9/aaBdqUtDJscarlnmcax3y/DatEgJZca7Ons1KeCdHQiVZ6PWW36GcD9dCyS1IsgJE7113VV
27wxnrYKpotmMbTCbpCihRM6Unwr4oKv9+9EuUsItEe4Jn6NFkjSekmv8gMb86QaNe0tOIZQXhsK
aR8Iuy2lZOSy97Sz0HTMrpGRWuCPtU4f28DLvNUAUG6TlKA6jDeZmAInp2gKZvzyUuKWkGH8iqpZ
miExrnsMPV53uG42+2XSDXOX8Mmbi7x81DipxwWgtcyT0Rq7I5jEM+r3x9i8noUmnT59igkK384s
nuUb+/Y1HNMqcMeaqEjh2VibC/fUzZ5W5BMS/D4DJM06nxB8QFTOL7ugIrGqVbUEOn1I8J3evxFd
PrDPmfDB7rrpU+XQZrgSSTd3Ce0aePT9pQ2urMd33I2c4Wl6FOW5nE/wsR/jqVZ6CJuLuWWyZ+8h
GihvBfa9gmxxbnfLwijNpY4jDQW09SRT1gSDaDkXaxwdtkbcxx6H7FNH4rPYnwcwIzDdflJ11Yj1
vUIPKhylN5uMbZGCyeVHX7vNUi2GVbgvhWrev1kQzOQm+DngnxkgJfaG48IekWh9bkne7uZKThgd
6sHXT5Ys6hYqbMJSK5bcOCsS3NzdmF+8O1bLFTtL1uzGR7PMJ6e+WXCmRBvbx2c72d8v7MHEC6NL
fdA1Gp3FdxKOzMdMmU2fOzty/KY3swqb1whPB1ODwgZfOXWpCGpChUYsMqIEzzhL33Ford0mmfCp
7exh0ickf/YWRFUwpgXKpRfvLdWgFbs5/2+TeX6xGGi8JP5oAO0OvUwibGZZcvKHg4SYkmv0xwkf
OlfqjKjh0BEDGfC0/A2auxbEivj7bVkjY5Pp6O1aq/DP4jCPD+6y5WkftahtUeIF6pieyoXhzO40
jACXvQdZsfl8mcZ5hSeqAZa/d6PzMATpfoXJXe8dqT68Bfi0QRdez7jvznX5R5plISv9bOuXVkSl
SPzGbPmifOmWhZWqGacXThQ2IG2cMb4ge9OZ9oYaqMGOkNhQv8f6UguH18SSFatO1e5CKOvBCoOM
tBTgup8LSU4FnyS0GNO6SAMUrz7uYDiuVbtddprTochCxlmhZ6mGQkRj4hk/7ddpUIAnhBBkm/fq
Od0gWbJ71XtwWZT328Y3Iw+4O7GmMx0ycdqRqmqRTyh+cPZY624415b5JSYyqfgWw9ZapuNPdLDz
tW2IDBFsTPVwCZ9Do5/R058igmGvxjF6O1pIym5tdq0gXZJqbYzGPmIeCBYrBHqpywz2Zglxe9q2
IZY5sSFOTiXmQa6N7Ynhh+Vo7oLZd6KNdEBQ3ebxLs0gGARfnk7uU4km02LJoapti8x5HVoTtcP4
hqLPGoRwrww2xLbRj08uRWx/mTguqVqi+lqmxcELsdBWwyzEYmkeoGqSkSlnKxhkoAPSoHNaMbUT
NkDxh57QO1TpX5f9xzfCCg9phWoxiLVsj0eBtbsDJMaG8yq+AgsaVvmIYkz8bYH1WjYYwh7KgCeZ
06X6/4GHYaB379c4CB8QXakF1nHzI9ErZeBYWRQD+ASxT+/ZXyzt81LHqkLeEWu6hxmaaLvNqJhQ
hGRGE3L9e3YH7BpQGCwQFatY7cDEuYlQ2T0Y5eB9orEeG00YVdGMgazJDYvpbb/Oyn9Bxuj6R1OV
x1X77DS90XXfyk8LCsablc11Hx63N0vEaU2sk+xblu/I7FuzCNdOoVfOfGqIF2dz5L9aNGEYQDJn
skBQdO1aWi5HzRmg4zzUFEi9NRY1xgLo/z8LC4Hu0nik1JXhT+RybzxRyCB2ahHeygKfqxrEEWaU
+YOVaTJIe+3/W2MpmSR1SaFQWnyOsUkcUavIbO1BXtlCFbsuU+ArmBCPdEHFJQcOAF7bixMP0nm2
0nlUlSE+t3yieq4fWP22D/4Ci4lqrQsieh5JJBdM/6NuQENbFKittV8mTnFf2YJjlevbsjucCDd+
1ur3fkcDYpHExaVqhahhlAQLOFzdVTJJM6bhvQImryOdtD6FhzKv2ds9QCRSScwEQwxGArPnrWAi
HkK3LKVnFkoL17bp2NWTwh6DDEoeD+SDknmh8Fy9w6OBuEynoJESE2MFOpV6ScBRkXrZblgpLrD0
UXLCngv2Rg3sVNiSv4FHL5vtlfGa1+t0Rid6xIhCqizPLC9p69ncHo/7hx0epFpslsht+0525Zhb
tvRo0D5rvPSraOV/lOd8zKSuONefQnlKra+w5O6ek6lH8REul9aOAEzn0cZNFs3Ejv4cC8hhIv48
vRKzlSPrI+mrNLejvY1lRU6NinoCIZRXNClZb0eapgbu1EN+cklUU5La6a+1Xu5D43ujwYcsSWBu
QdYg69kmnKsdG/CeJvIpZbqrt8esb5mMe+MZiR5u5CSAXiZdzAPczAmqFxSosvB9ffzTABIQDhlh
J7T5z2JroLbiOHyoQGla0OZ1OQ9pKeY7W732DNsYrumBWUbtIMYnmHpfUqRau3NSQQEyhdUIERrt
c25wwECvuljaIQ+tic6FSOgJiIB9pAds55fUUcD0Fa3nzNPYiEhQotiUprrddYXQcxOU/mlhLWTy
8FpPD0QuL+VHcDfB0SxpOv/orTRqVhl6dgjLq+AhnjqeR8MKbpM5rieivAr3GrCWZkQFQe74ajO6
VdBePwZUrxKTx8z0niy+gu0vcDd57v075Tjx9d0ir6eDm3nXy6fA21/Bc4AC7zTsaR0RBUEO0z3M
QalcXxS7i3iEy14hf8OoZQj2EjFQYFgjmkqo6lEDXHZLrp92XPjhIA7tsU0dTo1SDo6AjxRmQhY2
5/kGy25GvBL7K2xMpU73HmFuadVHuw/BRDp0FTQffsRvr81hB+dkVwqmTvSf0ZjBYZtT5A/zXKrU
cxsfeTv7napXZVWDaYZFw6K+UwI0zdXvPDj4WaxT/eH0Va9tOjGsSsQNrciU5ruaK9NkvwF6HXNV
ZnvRWdn5oc4ZDfLHiTORjtcz86FaUbGm018T8svgcepH1s/rcKZxRuFrAK0Azvp6m0AYAsYw8wom
MMWrIvrQrG3Du0Kx/hFCgmIw4fvQr8pPhZbmjxQqh/U1zYZLQDEq9qh4q6zp24N6uHWNbD4o+ahJ
g8EmNLojFvpkrwAE4dYVX/Cgl5Lh63xO24ux4L4KkKRFsbQrEzfgtQQou280I/I7BRt+ayzDl2q6
oSV2UaXeOSpfCx3w0tS7xbERuxAYY3xpMKAssZOW0+ASTj3HULv+sXP45r8WoZepQuf7+oPurNIr
iVQA32hORH+r2kJuQ3YCWtPCnvLPMafvAvZmfqoR2RJA10ns/rzUfSmJWnkZQqXTs1bz1Jr786Wc
zPQBaGE4gz/0iA3x6nadOdmbQGlUJko8zx6xhEDs3cuDp7xLCCAQG3RHUTFc3nuEPquQqfea7T/e
LQrNRJ/1tUARazhjwcWlnQloXVBEEg97SfQud4+YT2N7Ct8rJR586gryXiIZppUejD223Y17tLR7
w8D7g78sI7c9JToL7WGgFo6C4D9GXLdTia3s9PzZxxghhMF387PBLO/4BjhG9woXtMespFTPt2sv
cDmlDXl5vS3xiNIf1by34L5OkLXSMByfX4Mk6y9rZgNbTpX1WeDzMi9ZWenpmKksNZ0yhHoVvZMy
prvYzD8DqlT7PMDtV+UsUPxflbV/E2h2+UXrPjSB4HWbrPE3577cUjynqxJ6NFdJtvkha/emJyxb
GNnOpPjmMQqR9Bt4dk+ZqnCutM6ljutKpXmjPwiNb+3mIOf2qECSaNGgADp1WSXXkSZmLg6z+5G3
JALXaLFLi57GM8FAAbF14LhfDuD1dYFpbhFdeCBKLbFz/jgSlR/1sgO5oyhNUdR89Xy7CFWOgyWd
b0MYXtSmX14W+voT1JeaFde+EEd0u+MjlkLsRcrfmBJYDe3ZRAXNsTjfkfY/WJtuUmycaxoaIqhU
yTWmz786zNSfmOIiJdeg5s6MWU5TuYeScwIz8pHrX7dB4GRAnDL4xiO48RhPilUbjwncb2gKPDb5
pS0k1bJLHnTfFFm8Z1E3AHX6kIMsx9EcmI7AJ+VpVEQ+qFTV7FqumAKsDgF/41IkgX3TExMBvW2z
K9sIy6jbEuTeH9TK+hdqNjl3Wbe/agCg1So3xsdWPTQMCttprEYQVs7tvEjnXdSEtvnBAdjxKrzn
v6PBp4Rr7rr5R910bo/DrZ7FeIxQ2QrHezQKOwyNFivmJyFwZ2EAB+2fNM+6LvkAjTIqJwoSvfyK
FGMw0oN+EdOap5VypcKm/6xXZShCiI5dWsdkcEr7Y0AW4hnnIi3tb8blXVAfiH6XUznZnwUpaIkL
41tPubtereLjALveacKazj11ev6paqX3A6uknNNM+XBbt2UY7tIDR9jioZLFVC5/oqcvE5ylgobl
MIGwEcn0RiSEyi8qSZwz4KXnoWmkT1BKb++bJ4QEkEpMPDFHSjESYZ3Ys+ROzKCgYuPodgCXykyn
QpEVcJV1FDHaMif1SVhvXItdH3OKX6vZbm0Vty9BVjVh2iywnUNvn0DIZvaslQ0uFhO5FrJQM9Fv
smyRGZOY4QrlfjDwzvwxKPRkXq0YyYzvQZlHmDeEw9HTm7Zptv/huW0Psj0ipT7+DPUICbOtGEZd
URwjCelNDQfDaWlAOBlB1a9lz/qsIXrEmZsaG17fciqxixLDXBpL+0GUxRY6uHno6IDYUiqIxHmO
GXqR1fLBgy+olXokrt5Rv4hOnhbtHVg12dEB3ahSAe34LGOHptd4ecu7jiSP0t7PpX2WOpEdgL6M
KeV+w18I4Z82YwputtUYOZNZ0Cyb0w1Xi/sahsZlUwTKZ0Cc6XSt37UeYh+yxwNKboyvliMrQXhY
2H5jvND0iUlpeQd87VZaL9yNkn/a0madrDXyjzucmdTAkqEaGEKQmMX38Z/rD1tooVAcM7iw5xY0
Xfdw9tVw7vVWgTxhpLUhnsijRO8awkcSUhx4TInPDRrl7+RJIMSiM71KBahGQ7M6byOMAyZ20E0X
YD1lIxvrICZnqSWg7aqeUmJGAMb/4xc29lpjJZDxTo4h2KrHL0FbRHCV/xTuHtaTcsq3B4J9s+Rh
2ko35KIQNz8aOZVWN/qm+YjsOaMDaZKbua4aw+kerZj1slxxZnRZIwu+sazuy7lbWDrUzwYfc8zK
f4XmXibdidrA4XrrnA/tHpLISISA374FFALaoTQ1r+MeyDObyp2HM/AcYZOYzieu7rAhLlZ6tY3P
jNptz2Zusca2MveQOhuDfSqeK4VgUFigApJEy0LujkJYtWdJnIwF7NG4JewlxurGqr4tcDbmHYAe
vMc9MuiZLy+hoXMXqnuVc+0jCyMZhCgTWMrmaI7+AikXdgsCXSnC5pB5flWNraMKn5ylzqolmwO/
dXUR09J+PSNiy9VWL4Xs9EBIvIE1By8dT40NrW3vdMnCjCzWUhEzLcl+r2QwZoUN/MHMV7VwkK9i
vX8XOfC7A6kPUDBMY7TJd4mmX2pDuiv9kPCztjtjJMu1s8zl10aEV0nrqjf9QUtih+doau4E0O1/
xMjf8sBlYsQNAXwC612+dPaF7xVtgDPERWLXS26+e6X4wLAzLvPBbTE4K617JI4jl1s3o9DumQuM
EuJ0UglLc1ZhL4NQhgOr17rDcfjUEGgKvEZKlnB3QNvPJILIDiF8cdOUqOJ7cmOmhc2ow6hhPMa0
R2/l5v5L3B9Q1zXD+sF9/ADsiD8+K2bKwMB1SQJ33AISKWQ9jZJb2M/KXLPAu3GsEFpBLVTfpmGr
QtzIUsmbldRvOnxR7EJRvua605Bc1q1DLbg44523uFJy/Vo3iwZEyqafU3gwu6Z4SS6JSmhHTatf
sjXjtz2FodNgdGay6Ur6GB+ntk+oF6ffo9nQX6GAEZnFWOB++gKsLl/vQgFpg2pE/NTw2MxNCVOG
ngNjWFbyfRlohstaZ1DI2lDe7aDHk3aisTOS10EIQJibKJYYfJwCCn3Ykuikokm08uSmdcZ7itbW
DZ/5yDSleKqxRPOyAwLnHz6BW2ieOkINbl6gyfRzYHiXKYqGRyQXDUEwjFxDE5Rmun9o0ZZStvAj
+dE3ijG648YVlTqJV06Pwa94v0Z2psL7Ut04ruWgXeHgzObkG058/GzkKqkmD9ujQkEO93AKvEU5
/+ucdIJWUYdC6gixgw9cbed68B1r9V3619XxtzM7ormKi+DK9LgtNtgmnO+2GZmgRAB1JxKy4xYR
OJLoK4vhXk6mf467uvkfYIpxQwiqh/rXUVYhfCuU5dmTKTorHkw0oPdm9MB4NgTv+8van4omtmqI
oCFQg61OHAXIrGltZcBh9aog4XEu56GdidPjOeCKlrV0ljX4SgdExMh2les1wBi++p1oVC3mWGKQ
oJZ5IWtPYb5yNJXTGCotysRBAgxhR3xtiRZ/F6UrxLJlQlnOsyo6rlTN0lq0dV/pZeA4UIla6NYN
6voZfrA/BzgthlNVpCqBdTRuX2Td+tdFng5qYU2RlfE30HjfdB/7eOxAX2foVRnOEAo7vnSj04b7
cXqUT4GCaR+fSdrH5Oz2a1/bK1I9JyG/HISopFWPVgLrt/DHuqkDF9QUrcljXxUJoV5cX9P4zK9E
6w9Iv8Gv2ByLirT+z5fpqmyYRZsQd6qJ+kowpWyJGG8oKRZ7ItDIdnTpn4XN2a3OPO2FW1Z6k7Ut
zbzbuST5PTof1glXAea7Bt9Q/jc2u4acVkzcRihwyH6h1gyXWEL9KV6U1EE8Rpv0hnQDJyicrGTi
5p9/OsZWsu+bToyf+VxD/LUqvZ3Cc+fzhPPNL2E6yHTGqF5SWXaq3HjzWOokpVcxfWTA+mWhFn8R
oiK5++e6fi3bdPl9Ii8EO3s6GLzrW4plpCkm71Q5fPh6iYfVUeKlR13CXCzG/wT9Qidf+9PchJld
fXJ0j8HurmPy8TJkjgebKOiKLmPmAaxZ42KVwcx70c9LV0nTtxWoVWjzKqlJyzeDK+7VnUwiJJ44
z2s7NDdxvEiOQVaGcNLubxLgVLw8Ou5RPizRv3GZ1t1sccAq7OzbOZIbLPKItHS4atiK1a4RQHMc
QgSSFHjruDUFWJByP6rFb+Z/Xme4TYHyguD3ywaOLKgh08akZSUa5Cis6HtfsanUS6CBnWlAADHh
SLENaIYZz84zxZZ/ZRcm8HwhNl/gw0gNJ6MsD0iloaMHec+GKc2TtjuTdDXKrwRjkvgh1dMH0FGd
buwmutbBFMZ8aikBAc602r5UX0aRUb1L9vWsoixPJa9dWhKYDajyLbhtaE3CN8Nevqs5sX9fsnli
RrKLYuTD9gQ4nx8su1anBqCIpkAbp52FuZr/26yTDSLu9oThFxsgMPUJiDxO1m/jRZI6heMLy/rj
0Bq6GPFGKX5XktEvvMCgCXRX0in6wxHYMJTIH41fw1JExZ3MBEng326RzzCmNJIuyg0lVJMmmURg
fO10cM0DUeaVl5HCftJxDQRybFf2S3bcaNXHioOLoWW0j8+6lalnmRUxe2S7EISh+m6ykty/0fR4
j7WXBu+o5+ytrodgisRlVrXD80YwR6SpafIjiEf6lSSlOU2OoLLRDujfXq5sXLibV/iPBp7Y7QcA
soxs/eDTe1h8F4Fo8O/1uW+TY8hG16Y5lwtxtGKvIU25cHhIkyZgRpRML4OvEpdCcZvgyW6ih0XL
c8LMez2sLA7G7EN1UP+LTggnbT5EIxUkZxobQmixDmFCSJ9lfbvdaJPKOIcM9BDwr9Fg41plRYpD
KJbpaO3IyQPNkqeTYXGngU5zapPVg0wCAQOutH7FIjDONrNpnZp5+dbN/2e2fsyv9nMFZ9ALFxUn
5FMkX9NmPH6+57itdPROJJP9S1WaBH4714gBr0ubE4A0p+VDkiHDD9RwKXBWTz5tNMqJHfIgyzwA
34GzandcNXUoVXYqDnOex54fi5kWOTNYKTcq7csIHxijepcl92vrew0XXEOaG5qLueIxedS5iUSm
6ktIaCK1g8yuUK3E3wexs28Mfis+OAikUtfX7z2aEmY98d53ZKlhdKOKDb9tUneufvlrLK0cb1FD
UUnXmzdZJQ9c2AQa6UnifkB52YhzLSw7syeaZkkl/5hT/JvRaAXZcOGqgDhxu0Ss2uhCJ4Qz8pJq
SabqC585myer8E+ojV6GM06RdwdNFdDMFA+80CcO7o1OhIgXSLWbQc+uawhLvYWcALmoy70hiD2U
YEftRWWpPJB8Edy3pco+weWnIngC4r4D3drhj8tWISxebzDo4v0/FnJ9P6X+cy4B1CqqBksKT1Oz
ub/hhSvsVa3ihMvkHv5+dDC+Lxbc3aM5W5rHMFvHhHst04KtJfrwKZKcKwiWw6VBUiRY/fx1DB6B
1c9PRe1Zcd6PVw6h5rr0wHKIjz6UptLPkWg/qJpmPupzvrkdai0cZmE+7uggMVOIBjztg5ucPI8Y
FHauxwWZ/lfOTuQO+WO71IS29nZTKK3ij0qZJJX3lAT1RAfCHboIUCTq5gx750v72HuHXMaS87M6
09jnNWbOBmEj2/Z3DeIIcEVj3d3DSD/No3fSfEVwxXFZo8uDqqX9VuVnxOYyh10y8Yan52Kcmrot
cbibUz6UVhHeOvX3XGa0ZfkAlUyDyRxzxwD4dcv0RGrGGYjfkd1TGFV3qCWGcij8DBNFHAW/EEWN
vCehxVuXwlrbISml/1+9sVSV7O7JYlr6j1wrNWS0+9j043xoEi/ExwWG03+nfPIxMf3q9xi+5q11
kP8/KVoEyNfy27zXRbVh+1YxOAQwI75WjjJumkAZkaR0TNe2HaGLEVyamJqpIORyM7oparr91O4E
KQ/hA1p3YZ9SBQlZc3Dllts3u0EmQnFVjpDnx2oN4ta0K5/32jzYclsJdxaLYmzF2fTxkaMwWsMe
KJTQ5yir0lgTd5OGd+cmKAhdT1UpLlg0M2dOZOloR8BGQ77iCb9Q0Gpl95VbgZXCVt2/4A2Maxnp
vr5qHOV5SqU3ap10Z88dAuQ2HxDNC4I/g5WlQR7ad9n0/4v8xYXnTHVxQCDTC5zUYW3kXdvbmAyw
u4KkHvS8kOd1/UoLX/JnTdklM4SDliuGYmSC+4DPjk7P0kkheEQ5bvPDzeu0r8A3vYW5eh3n6B8x
D1k/oUM0ckc9z+RDL/F4GLosUDPzDqZAcvAMYDW+A1QGo89s8kNik5i7n627xGOcqoKFTH2VKjS4
bID1h7tv2JRBss/inymAoGonuvZItNGBS0pNBAXzhhmYvCT81+3pRRo1Suxm5Z5k2P5b6LqeanFV
OcgYkbkqeb7CM1szfTAGmik+b350EQSh44Uo688+R3kMSVIpBqU0is67oxIpMA1ZEkRPq86/vodI
uXe191XQfldt3mO31bcG1JP/u+73jDhpCNh7bifbji9OMRZrEhXXnOqexS8My72TF4jBZtrWD5Y8
+2vSu8QgfrEg8422s5AeIwVTgN1YMz6M/OC8JnI4EstlzIoAok4XglpJHFgGWIQJVKWaanuyxue9
xgJz6Ed7mOl6mVlEM0d4QfB1QW6t+c6QUqXW68avPQMPOfbw9aBhNbE/sxS7wTytzNF/tAXqATed
LsUKTW0Okm7eIt2XatGV/bcRVjHuP3ovtE0PISjR1GUA0bqRHCpbB8cc1PhiKWeLrALbB8uBbDjN
RhiyKutbBDQ5BV3ew8lrymleXI3JcbdshGiTXTu1D1yyjxvhRXaKoDmMZQ7sklXu+do/eSgUWRBU
lwB0iSklucQl7XHdPGDIM+4kk0CdvfuLfQvFsnXWATS12ZmhhYgJ/hdWF9yOC8Y8p1BIMpmOGIEA
oSMBLIP6glaYann9o1wLKsz1W3Oiz0slzhIrOO0yZhpFbSXH+9J7YrVJS9HO79LUgofqrAdYpzFn
JtRaSA2VgXtdG3uXx1RXvk7pSbBSalxDkjipi6tuohSUY/28DnFmeQrvYSWMWexL4IACnB6/skAC
QaOcQvFJ5koKcOO2LJDXAWqMCgGWgmKyqn1kWuMQKphNSJPACJFJENY/aqPcMYId9XVjCK09Vju2
mCmD03mVs0jyBROluB0DQX1ZPg88/h64Fa7NHuMYh61tvPyIa8ER64HGm6FI6WbrRQGTupflyw7t
ZlWSfdVK9cd2/PQdcRgqOQ6n23mmH4Ep6NmUcCGqlYljoahfHOYlEq0+2qse4miD9CiguuNn7Vra
W8RiApgBkIkbu38yC1qbFmhLwkpGBtv1O6Fr5tamKpZCotb/vbsqjYdCE8HykbNeqhQV1uSU4opp
xc02YjhBWgbSWaHxK8pHWCj2LPn1Jd0Loe3jx3j2BxX+lYZS4S6w8tpo6TTCkNS6YZXzBrZmkY74
IyZSXr3VudQTgjYho6gYmSPEj+r6B6PPvZXzEmi7hmWS0f81TgMbSDTITusC2KUykWY6Z6AOKvKb
SlUoHxRdNRCooj0SHR1SCwiXMVhc9EZ7ub/CL+nI34qaqUhY2jJb0OEd43Q2MCbRKLjnOQtUzEis
kwwxRsFOShnB4jn/21ni0fv2mCZ6/BEKyZTWrG+Ioff6uOVZW8EcHMma89spG+KiFniXPL1fe02j
gGLzjwLupqXpHAjjqSnf9hBWTRLMlsfgkHh3xTKmC61EjxbElUVtUy4j8W0mWsaRT9kodFME2ci+
F6xdn3sjV+CmYRtZZ6J4CL6Sv4VDLbKkHJ6bfSPCOWr5txQw+xv0EeIkrBmCLYwSUikLbIxefBx3
ncbq745bGN0M3WDveA9LFL2hiiStf6P88JPzzSDn9TIzJ/ozVLp1G0p2I4rBTNscYe7Y0/ZBf7qG
Joa9J4aOHwWYl8LRRESXAk1sJeik6REQpe6PJJsPKuTO/5c4fgSI0or8R9s4qAQ+/bKsY+Q4jsd2
wH7uWXeUVebsbuiT1O1o2oMK6Y7q28QTw68V7boqHNk+AEjFCFO27ZBTifte7X4Wv18VmZ9tdTOr
bGepeSffGdvY11lzJ/FDpKyDECsojih7nXIXcJ/f4oryp+3X7aGJxDi+ltURUfLxPonZy5w4iDf4
rzMTcTkS84sE1ggKzKI1zr7YqK10MvKMwycwh5fdZcc+2T1yHBmW9GEcxEsu2HgD9S4m4jEyVp8z
2qqLB2xfm3X8QuxAR6I7iYuv8HwOiYZFSsot+ZlmDiC5XlVrSun0W0Dd/QIhIdavAn6gQrQD+/6N
3G5Pg1kjJGQwboSPC3Y1xJqK9ZlRkoU5GeA3Lm53w2MTkPtW/h5Flxq5xZq9SyF+EDXV5EhAG89y
AHD4lcPh1aCRQALpZ0WPKxkFSJBTz12ia9PMqp0zw4Qaj94MRNRUxdgoE+TBkrHdV64aH93Rx/Lm
mBCWia1azg6p9htVjhIn/KUZKfixsJOB4npB0ZpJ2yvgxcDrLEp7NXW2VF5H2eeFUyYlnmOzZqQf
Pl1GVzyf3gvY6cG2k4RDj54uuqgbBVthZPeaSGO25TYfD7hLhHK7Li7pH6vD4ztPZCqyX96PQu0c
cAXUgdSeq+6mxBZlnG86edEPe41533UwRo93WbxW8u9F3wNHYnLQZt7yBuy2RU+MVkYiylGxe4X/
5NSvlhsurM+W+gvDAJU7aVKGBRJkwW8bdV7ZM7K+gH7oFyk533LEi+taqHbTx98LfSQSpCcyWVEz
pXC28jEJVgz7zYE6j3lUnnFCR440IxCbG/NvsVFUPJKt8oaspn+Z0GO1nwaXcEmUwpNgYXZn+OJp
PeCqxWMz9evo9Q5AFa1QSbE8/L6OmvCXJjyYV/zx5InJiupC/HkaZXFIbF5XWElpFeN1GWEVFbMt
H76Pk/PNq0SYvet+7ktmCbMiGxUEAYxC80jYPk5XR1gMyizuRe9hSJDEQh3mH0iqOOsbmXbz+czZ
c9YaJVpIgwJMEf993rCTzHcunSEm6gm75BS/l1+Xg0X2SrHuv7SUfA1iDe0Mm0p8ZwgbuYIGccii
i7n2jl6dyes+vLCehVWb0fwMmTbt4VTOMDtgV5MSiqh1zdBCUYHYPc+CaTsK+MrH6uytbQJb3O9H
lZkaQVwCh7xJRscVM+mA+SVV/cZLS7fg65xM5rMJYvPcPlOb5oXuzh+9iVSLb4oqdlMBrC+NavrZ
2vEJb0oJE8R+nZCb5mvV0tT0S3g6vkHBjYV4x6HFkHEPZSQk9iiBWioqYLdokn7Gv8riH1CRBkIp
f8fr+CQ3O+QhwTZML/PNgGtFWH+8tJCqzTU1MX3nUBPFeggzsXXEQsmz8C4Tf0L0irs+75mv2x0m
BP+jrVIFdr7stFW8LielZej+UzdhwwDnOxx+PL5Uhr2L9g41pU9QKfC3BysiVOMGuR4vN8oG+sHZ
DVA1cN2nPGobW2F6fv1vbBaghZ2yO+9dyczAIG3YtHBo90x85DPc15JBu7dcBGnW0QHiclTwWqgJ
N7w0yfdmaF0JDaR8Kqw6AcqCvWSc2xfiXQ9yL1g//YhkKnGnEqthRPAapbXMhgVX74ndu7D02oYa
j3IOEvipcL3PhoH+Klf+TlTzntzHdSalVL8fHyw6keiU5tuppiTEioPEHJN6qMOdMsF3l4HmohTJ
PFrCHdbYMV/icUtyxtp4IGrCgXmLMvQh2wBnOP9UmYKh30NJNNKVPR72qxawra+AJgIaIPMRdt74
iUVCsB6Ei9AjR+kwe5xLt/CD4JB5senxBG40woY+/AmzMxr/ufuprDxEOhvXzYiniINGPqmzw1wH
OFunm9ko/TdT5yWypH1YDM3x3CNLdqbJFZve3cgz/r+NLslwV5fqKMrnA7CXac038Rls/yYNFv9p
ahA9XAMJRF5VPrAbXgZB+oAZjify98RvwXiVP2MQkab5wf4xFkUf1Oh9gHCiWiqzEaWA0AvbHI+F
KIZshH8Xd0BQGZM5c/YC2SXb5z4rEAO3lw0xxqnammksUuwZNPPfitlcmKIQqv5Ap9U0VyBwtNUp
Qvyr7eVqcI6lW2dXELdt3yPxUMoD5ZzrZFlR2ZleU8n6nugIGZwxJqyBmMCHBM304TpcpdODSIHf
chFb8eoX3JMX8uGYfOn9k0Q7r8SpdZb3EC+SKAG5ad72trYSO4gzqLFpIcgFMO5zI5vVT/7dPMkU
OZfxTGH9hoKjnhCYnMUf3CkLDGkMJVSZ7zyHOYqkoG/GKYblsu5i3mEjzLWyeszLma39uiSy15Gf
gZaDDuu9ibK8HJUTwcf4+KvTjkLrRzfB4ZzVFhV7s3RbixWPVGb7Nj4hcUMy19kLtnOtGVZgi0Ox
9D6frzkOF+sKFdHEwE+SRl2H4xWMJnHxw6+HgkY+YJi0oEnEcTMBbxLNhpVruhJaqkjw1PmJFJHM
n5KvxCbuKLFnTL5W8jxLbrwMpU0dRPCOsR0Qb68u9FJqDZron7EI9S82Po1J3VT1zXzRVncLTVGo
52ALHzbDOHUM+YL7vcX05An+k5J1NnaTr1Ea+czPS+YNsK8q/wM+B8MQpfoC/mOEtreovNTBG97T
hT7G9jVEQ/5SPV+bjkH2jK10Fxirv1zra+CJFOV1MwnXvB2EHo9I3FHL3O24MuchUlfe5HgJLjlE
x0i/edbYCOpmGEhA8xv1KrMtxpQDpf0+9J4Z5VPWgqhGl5UoIyGXU4+cF/u1gXW3GN95CdVECVIF
IQvK9rJeUayIH+9B0m+8KccovNbLoHM42+drYKizJExwkVce31tM0i+Rk7wIJ8Wlqe0wTH+orXdN
b/upPardWaUoC4+XTVFPBOhJnRor2t7dmWtR62DOaPGVfhtpTkqx5JQlNAHgN451Q6x5gQrb3DkR
uiak5K4DXFLzBiC9RaF1q7pJmb23GVn37+1+QSMqL5p+aflkf8FIYTUoeC6wCLl/V5gHCx4wtxe0
uTN3LL5WBPYlCJ3JRUM30/LHWdIf+vhUI5XCkase2AFBKXpzqmerm71sR0BDLXJdEN0YWzojkiRe
DDiXaAUZGJR5nskmi9rctCD1D8kRYO6OOVvoSKS+Hifn+wLgNQqIAIOzTk8EhxxKG2SZv9xKFob1
AkxIGHWezP0OipEA3y9ux10Lr6hlHqLkOd6/Sc9sO9EZ08eHuKNQeOk4ql+x31bvSRE3HhiqKlmO
mbmuiRu6DrwLyUuK6L5ihBEHXCookTVrUWMVj/uL11HDMH22wPA6NJwxJNJchpI8N/6K2G9N4M9f
l3Fqrezy8bjpdVcSKP0j+KVlVtgA2ed8YBXTIJb3pCL1AoYSCpTpVa1cZ2eSSXyrCWI74fYNbt9L
epOolZpoh483025a/pi8hnhyOG9Jr1QCM5gaZMfG4aQ/wH0HSfyRQoUKXcbRvqgNqc4IZHEuSpF5
r6Eqn9Kk4F1IIEQS38ZjS9jJgQOnY9xi4CXGidsNF/HL8+oiCElTYcM054LRENxRXf6SgAhHgsyE
XPaxMxhV1wnL0hwWiQFpB86uM29SVDxUoFA3ZFrlWczVyaqGf8w+Q8X967Jfst8bs6CdPqdyy9Ez
j15FejJ/RkfMTEynUmwhWAu8yn+rWsv8qdZ8Dyij4Ez7zDGKjOdtwEdgkWp+wresHjwMcqWjfslR
CkOP2/hRcnVCbOk5C82bFROCcfVY7BavJzvreArgINRQFjYrz52DAv4SCoijlLoP0uLTHQiz+ulB
OLLxDLUBmzOkL1omAitA9xVtaWZMZOBZjwHyiemKD9SBPPgb1/sgTIHyjm8oLRS1uqthr1SKL7YE
ZNeiUMdGO4bzRh+M33P4AwTayK+9GrIwFYUe0U7C3Eepgsq1O4dgbnu2GxP4+9bRMZi6fbRgnJ8O
SA5YSBHuMAsQq6yXyd/kHF/PtkZvN9AI4ZhMKPIWj08Ot+TMFZloSWY84eTj+ZmuF49CSL+AlF/a
lCyazr50WyxONfiXh0R7kIEE3Kzsz3WhCflsXxJjtdDaEh6dIA5x8GIwkBQQrW9OzXUswIKvrzrc
3t1DTpCP2oPaQbK1dOQw0v8b89XrK2uyW0+N92JHNs2tUi0JeaplZ4Xks1pj1ZI+V4oFB93Npqjm
noZdy3kOkMJyHYs9EbGgpf9qF2ujNWjam9JUm+DvppP5Ekc05biYrtpEDLNY0SvdvvS9B75LCPX7
3qYy+cawOlSoc+Qy/M5o1p5VdHpSbDJGOKgqcVwayCwCm9iOD/ri4OM3jopNAQMRuK+CP64HR4Vt
G/ykEjj84UEN8v0YVVTWMxpM4Rk8u2cR3wsAujpKZ1mbzg7iyvrFFGKLr8SCf2ni3kVUv+bd+6Z7
h8VFbh2Jx91c9VbG0DhAp9aooJZaHL4lCSP8YHhKyyEyXLtw9lN0VZIR4p0+zRcQFucgNwtFvtvK
p0SGew8QFUlttDk7lOAzBbCzO3jLX9K8hDwaueefT6cJnOe3/35jGmNILR0dv0iVvWF4EXoRyypx
GrUx1hfFz+nQevCW8HMPXywcef579NygYdqAlfiCMiPAZnMI7pF62wHpBjyXqiQ9M4Ehz/fSXImK
ZX9zwSOmlrRYxixeJVhe8IL6gQ6igbsnlJBfJZn0BlOJi/z508EQIyswZ0wU8ckVP8l0X4X+0mNi
bZX2ssA+4wr5A5EWUppmPw4ZwdtcJuTjXmbfqpA2/O42Cp2OckiUw1a/EMTocdUMb6LMFOC6vE53
4klTSY+oCFJf8oKbthncQtWokWc5nm7yHoeo0XrriygGk5RjnfXiX6dGYOpZFfba70VExZJJ2gez
EszLVDtvSElC1c49cEulrPj5O2ZoUWWjgXbTsb9etV2WaVIVyE3Qquvf4R5jQz26JchfCDHDLlMv
rFXNmEY1z+ALjFFaF9htIPdy0NOeprccnnE/HCyimhfqG3VkeGA58CdVcw6H9w2o9jEaI9rZlfIX
T4g3ZEPDb2ZJDOk28R7HnNH8s9QvK9AUZ6COqh7SPEqVqIBbybL7mHYI6HmOOVZJsWXvBZeuqDHF
+JRVDsZHSQic/neL/zxDDRNiljG2nMC8nPRY1c8Nx7A662YACxblh83E0dSt7cjQWSX0ex0H/iBH
yDV05Vr76TBQ6eu0w0Y5zBf5lC7IKlZ0LYk3LDTgcqCTUfGXugToPrCpU+BqpVzgvNflxrfBYWEQ
NiSpMhIP6tg3i9V96WRo85f5GMQPa0mJaEyyEY9RwfBIIjEUq6vF/mAZaEHG5Tk1Uvx9R2UGwwx/
4Ax+TLRiVDgI3v9104jOvZ3MVNfVHG6mPnqjBp+z2ulZV21RhKpguH8QyKocuDdoq33p3DxGfZ4b
hR874V8DWGpF+827LJ19OHb9OZ/OPPmlme4rQTExo7i5GUPhwpxMEeCQZZjUvON5W7GN5+SptxkA
H74+ovMgNq9fYRl9UQXbnEVm5lNLuUFCoY706X/U7oIFUPVt43YSdTPm5D/TduxJSnmVUmetm/Bj
TYBVS75/vkru8HpsXY9NuBF6M4rOznJqN1DQaSQFqybabghojUkC/CoF+gcCNMyULbSHVAii961v
/OEhJY+dVJEBT6Z1Bvmvkag5sGWD0Ov/E8dJB2LSRxHcMPbdWJbBwaM2dr7rdCnuJcMD7fZ2Rieh
byrenAZyCVuHfe36vGST0j7OLwrhiYUSrDvCHFIk94ze15X8IE8/YW3ZR7OO9j4LQnRUZr/T6anq
pi/rJWkMc8gql2wFC9myaiyv7QO62eQOySfoHn40ds/dB0IyayevI2DtubB+XvYg9WBUHobtqNIW
1XP70piyfBgTyAwA3p1F1WCDNlvcaHiKxch14mMph2q04iypCdTZvMmcghr4ljuKjiJjhGpoE0ja
ccnwGOybnAEILb18jgvLTTkYD9wJ3qanADbKTcQ3zUCiqsM21K1ukjPPBYmvzlwLIfJUxorISxV3
d3D4KEvV8jCQetNfTHRWiyE5qV+x9jtQfSFbTA9vrR+Xgy0pfEoxjcQ/2bhFcKSIVL526qehBlxt
f3a0CUhUtky4NAC4idAtGPZsmCY0y6BXNtEc5LfRsSMZyOlzRtzOCFiqrfmHOu6zAL0KXaCIJ1kk
gI+j6FhaM2ilOkWI66G5GaCi4PxVkTy37nDwaH+jG8TfRMLsdODEJVoAt1mPVoqoxbXFDO1MGTtz
ctiPiw61YuEAL8YOZCID1I35KziejmXmU2cGAKCM6o8NGHYv9mgr+AEAVHbcZtYL3TKjMqrn67Dc
Z29maIU+vqMozKQ/OwKvFxUqxLoYbMkzem+4uPAqcxc+0rAsKFWIcKX+mJ4GYZ6RMAwXNs6asOrY
r1YiX+S6EgihIkSZF6krJaphmuTO+TcPG+jHwgSmuqvOOwhOHG8v/BgYY1tK4cXa8bw6nDv0NpMZ
NB4RyfTUGm7l3gGcmS1ug0tHNtMNXFL+KqAO4H9ypGN+IttGUb9oRGH/b711SwCvZga4Um9G754a
l/adcOLKeu0qswu9wu08l1n91PdHWKySoxja2H+hboEIbCeHuSY9moow1wO5Jbraj6LX8MoygOCX
EG7LpcUYfJ9139iV3AbpMvLs9m1DulGVKo/ygIhiFd3mDvsBp1DX9/HJIZK4j/UU8ptLJ5f4PADX
u5sH2B1Q1QdHPfO4munUfhmKpnSnQnGNJqwCtC5s3yuWHDIely9okIlZujPgejQTKiFnMGY+1Cmt
J6syXLuAOSGohWfw53yEJjyb35xKVkQLqZ0A4jqXJVMK1HNMLOaCZwcXwaSmb6CrcxbU98c28kha
BWbKmILMMz2P5boRDCC+nEMgkX9GADU6AMDGCgpbJBP8DUMn3maTEbO9FiSBPX/Sv73cjDuSG8sP
kMNIZIIHm3J2p5YFsqBtU+WeQkYZ42j9Yl4me1KZUGfCROlL2Zfikw7fyi7zth/MlmFeXL9+TA4a
g4mWAAw3GL6+ctpiUEpcwr05y4Uz2o9U86w5XoT+u8pNWn/I7r7qCjD6nOiw9aMbdRgvCZ8aH9d6
vtX31ylNSP9NdUP49UY9SB1bIwxNHba5jj9L6wVeJOq0fL5EkQKaQpSmMNRV1BURFst2eBFiIkqa
mwsIsxW9mUr7HXLNmWGujKHVwphHYPYo5r9P/c+2c1pEvp4uTN43uPN8wGa0UDUAbaBmy5gA0ohf
R//W1GlXqz826KX67SGSDd2aG2IWizvTFQQtT35HhBNcTZ6xG0yEeef99a/bHg2cqv1qYhS5aRvh
pCTqdxuR6/dl+yV9jjKkbMudkhCNQUA2EdHJtWV5mVmPjTKXxtPgak/ObxI1W7thTaTeNKAhTdys
X3U/vd3SAW+D2KXPyIb1KYAXietn/vJfT4of7hvLGHFxBBb/TSswFDjm45z20jII9mpUYdYyUuRr
qoosFseKRsttKPMEaAiGBqSnPez176mSjNSMqLZkQtXMfAVuWqhK+HVjVA650ixEbkCqJPcxoOWz
93irIMGbeAEFDOGBz0QR/wGpAXvrt7IRvMZW2QWzmCilLD03qjlHbrU7xraxAr3K+l6WD/1gEnz/
KCn9bmSeUaYahWRiTq/qZBV4IwddQLcmDfMv4f01GM4EZLlyd6B7ToeizEsZMI8jsbAYT1zcmRRS
giLT1balqhfo/j1g5FfThvpTVmIv0RW72cIekYvvjIK7qqMkTSKEiopLdwb6kM8SHzKO9PY711C1
riH8X0xeeGs0MCUeF1RaHsIdyl2zbJw8ppydGhLoKU38YL/GXVaECjK/ORQ2yWVvic2BvxNItbrb
PRk6HQszbEaYoivM2BX3IWlSYbqlp5OqJpqjAsG2/43k4IwdnAB0sQjEnHfaRmBlQHpi/utuhAgC
28nmdh1BwkegaTaKGm76/QxIU4CkjH1RzL7WHFagH1gND9YUgazuBdReHnrpsrOOaBO0cZ26mWaF
JF+KjIb6X/FDwo4uNK1Kxj0pwtRPpK4WddlM+02cdxWOzjmzhylNf+r5RvSI3e8J8NbhpnQMRuAH
mwwem6yeI0PXaQOftb6gKn6ALE8P/VvNFA1FrI+1qbea3bIgTG5RKjzPuCQJ7oid7mVe5lzqgjm9
eUi91hxiPgY+OsQskUXpejcPywifxsIzcIgMCjT3fRp7N/OhoA4myQMA1Ea50i6l3sE6P6yP+j1Y
ykuK37SzaQxwiIOxwHja/HHLF6wYI9ofNl/DBAMEO9Dp47px3mjZ0geM9IUb4EAagHZeEZYiJ4qJ
3WI/TqBhC096DNss9MttYRZcBj9CDwYJN9mj9BBeFXSiVeOhXKAsQakZgrl9Evm4UEjtXssLI8GI
1B0fBIhlz1VkQX3NTfn+YR78SUWmVgrEH9Zugq67GnJgce0MxKHgLRBM1TaBTI/1tKi0pvlcXmXW
UTqUJyk4ZfuAoJFfQ/2xqfYF+7su/BXpnzLp0GH1dt2DJIX15AF4XJCbA3lmfzsIcSP0I83Unqf7
IG+XvT9d6fDwPn8iO4TVg+pJ/mULTh+28xm1shM+chdCubz+R34LVMXF+GSvXGQcfeQymOT0EujR
wscLv8W73fhHPejwN4ZhtBNwL6NcNe/uvRR8DB41nh/8YWOlaWY5tYgI0tqg10Ei1DpG9BGsLVIo
IFJjh9wcyF1TzU3c94JNikcR5Y1d3+yvYaaVPhK2/hwxUULL0JZLToOG0olRYuZI7RupRu9mVbjB
Q7exLrHz40qJAuNw/BhGzmvzflrTHx9Tsq5QI67lkfs5ulcUhW6l5CHCQoiJmPDMiiECyAYVisBS
vfDidHd/+CA1cOCEkMYLmDw2+yeX9U0rBFqK8UOgYGxvNDXNLrWqc5f+R5EzUriKzO1NX8JG+CAS
ZjDfO9bGefPE3Q76DjZSbMQFik/rWOOCJNUFzG9k9viXBVW4QoMZbG+W5aT0V9rKf6+9lR7VubuL
8XsXdeyBzOgSdux6o7W4xmMV3x0JhJFBy+e3WFVt54ULrrwO+Bbk7GVj5LVoxT0ocEYzHkYXfbcX
xglBXkgxcdb4ZCYsbq8iODfUj+FgX1EECWOJM3KoHJ5OOizxUonVZezwt3+cKhHP2WDbnlllqsZS
XX1nics4EvKR3uee7/y4VQoLVHR58LVZWOYH+EcK72sRZZWpvYErt3IbmYKgJUfGg5Luf9iHHXpi
Dd9v9wsrmqp48odgVCRtlKuECt2fA3lrGC+nO9OZsO1TzOVbTYQubLTegiGu4/Q/fUZYKb1YALgy
Z4MOoWre9v1ZGckasUaybJtJmTryuE3cZ9ISCRWxdvVQj6+gnN5tkc41nSICHUmQBCjqCp4LLPL6
kRaWFvtQwAgEuX5kvdHrU5Z3YRPwg9wuGp4pcLY+JH+e6QX9M9r6M7DEJX9pbb/9UmVA1GXKanlD
R+1ckUwBio9iEygk9zAy42rWK2T906NksI5tI1P3JvGiwFPjfh7h46wfxUC7P+lQnEXi8BEIxn6U
/aA/25Yf+pN75Fujb16wG7HmJs7sQZvqHAHoIyVpV6Beo/lJ5LkQDKXMYzKc24XoI4QdP/LZULnN
+yWPvNCQoJlPrnSxsiqVnwbiWZMthBl3UoZrjxOV/KFKA9nE4ASfuEtYX80OtZJJ8kD/p7JuCcsA
ANhmszxnm4dP/3cym6xl53uUBpX5f8jQOl71F6N2hGlLw5ehlt/ZUSymGXXP8dg0iBMqZD0bWC2A
/jUlUhWRImx7O9O9mEKES7mCUyfhMAbBDFH5PfgRDYEMnZHG/HhpAeWR5RobZMOgrPD+GdEL92ew
vH4SX+f8dH/gIF4Wa7cZlHWf7Mle2D9munZxwy/bszpoi9f/mNfBfHUj7s1adJxIqut7S1vfYKUR
n0e1/c/JsWi+W+YPxUMJj+8GmsNTSpTsulDF5gto8avqx5E1jk2xGFCwiq8Rc00uqh0HcEWYfwz9
3fWR/qPMs/KwAzd6P0hHLM8DJruEO7B8nuzlK21Y6WWyQtF4kswufnOFDsYD3vgghUgN8YBQnath
WNhoPK5w7z/wJ5VJXePAwJKFEnznnLq2FP2YLtk5ivGzoO8OzYqIS5vB5UOynbN8f5SC7ncNAPPU
mMS2+eRp2KWrDN0IDZLZsJgoDPyOqjfAXpX4b9qDfTfCgFKpslCFNQ6+He3T1GF2r2YFOZ1TorZc
C11kg2tIeKwIhVL+0y3SfBnqPlzsGJIKmE2+OjPf2IbI+JETKUVWKKsheCF5w3Hbt1zPgQaRAQhq
3l+uGfbB3jpD3XAVVFlzMsqKKdbmX6qGGvkDIS4yh8ssOjAvFiyzwIfEl9GZ3SVCyLrrgg5CSEem
bQd3RGzhP+WYwl4dz0U1vjj9nqvvLbKZmrIBwDxCxjsO0Y2gTBM/svVYyiQYnPT2T2oOWBXByLJ3
cWkdjnAk3opaANIuylvvrxaVtQaN5XkxYesLhC7AeewIEionwno9axBtkNiCeTZBYRtmyC3ycG6W
U07UcNzq1huWAMwWF30yGQkzVvTkeWw9tmT4BxSMmDYu9oz2rhQCp/1sQfsrO2ZiXC57BMYo//3k
JcMOFPl7Bc2K+7NVgmMBwAKqWTY7Sjp8vmuc0Rae/zsDP2Pkb37ikfte0zTXgtBuSVuhbXrOVt+5
waiwWHqIEgpgKfmJt+57/IWETmXfhU/z8khwcRMX/qwnCQYvFYvL7TzMmXA4iu3+z/UVm5IF1HiJ
bgfB2p4/xn7qMK4ZWWL8XDcURBqRK4vRIpuV9x2ECHr5Ytn9kvJYpam17ILMXddWODruTOFmMNkp
bgFJwjhq1le7Ghm8Crn+VQqGTgzj409ID/mJrqH2rVTmtkr/VlGyYr1BpZLOUeaZSD/KtPR/NhEa
miOHPkwA8WeTASd5r7E1LMhYv9p6v4pv5BcEsrJpoVms/rRLBBfSb4A5pI+UT1hPkBr+hzFX/zW8
Vy9dokQSi8pvIMybtoYJF7ZkAaNPiRlOVaq810aCh1CdZ/HEa/Q4vfut+nxe44zgBq4NAttvEAon
F2ePnIO2PkOXXMlz7vOUbKbz+IJALoXOCg4MWw+guXLcl8M6F4sX/FiYCdRw4titiCzv/DM3MuLB
nBT+RQV/z2Gg2o/+O+lTw5m0H2NhzJQ0XExsoLTY+sEvtE3xb8cEjW1oPGszdHnEC3ZyVPpvmB+Z
inxhBYiltpv9aEgJh2hhcWFXZv8aykL6PWaa9jPUEsnphKc8Gn7vPv9SHAuNz9h50Rfv8xfJrigb
yl06iJ1mQGe6x6jv481EoZnWDq3H1i9HX548+xFt27ch7/vJM8V0PEHh7DUUStBaPv44SLmkUYwD
jaOAhzWfI3XKGerOJdhHS0A4u8CrFHWR3KbCl4afEtLhe/GchDdgn212WEpWUsveSVs7erHBKPKH
bwqAquSQF5nyA35gNpXKzhYYWzAd1VWF/dJRQKKYXt2lUZmAMb7rB+BY9UXec4n7rMjrDH0jnp7v
6FcUQMQb15G8X8aJYjRSB6SrNlGxLqJckVTg5XYQjIyqctn8q1hFg10LYU0IWu6OfvdynhdffqWN
PgRrLCcTQVMqaQKfhZ8uEH9BqzoJlgnm775n18ZyCZGNSuUeJEA2LGcTsBSp5ElW85cVJH6DghkI
WfCVL2uKp+rR2QMK+waQNKoVVA8vymHiLRvkAd6wcnextXtoAsvnprr8Qe9Zb44uSvXD1+MmlYmV
s9m5qBXsBweYzuooVkdb2aULxpgsrQupsCV1sNhXU6BcqeehwaWn0IA7hwKd9z/37Mwyr+179NrD
MhYBD94tAj1eg7ug8s/KjNkBsOo3KM+TIUOa+IKh4fmuoTv7HzaM/57WW0487+4dh9CDH+RM5koo
tphxdz88kvp+v2asGWEXVvI3ySlxx3HhvHjadoa3aP1YrApfJJ4cRR5jcBz9/7ov8PDkXkOvu7m1
K4dSBs1uzAcdBEHFfbYaLBx8bD1T8BiQl3C06JD+vJ7/sGuDfXFRzAP3kw2TMlBgpuVdgNbGyvrg
R5Lf1d1M7Zq0meqDAg9Uo05cclk8I5nskphUtjVAh2Oszd94kvPAdXIpxVTp+CPLnsgRIYXfq3Kh
vMfSIRxGL+VMf/gLFGeuhqMieFWbIuWJoCSzdfou6xGZswggGHZ4y609zZ2u3j6sPGwJtEo7IpeI
tjxd/8eT6DxYU/ryAwYIlfP0qK54ypmmu9doPc7rP+IS4Hj6KMu/w1BqbReouvWadU07J0GlMXHL
/EydBZUVEzgSAM+ogLl/yhlPliKKs2R2Mx/gZMyJBGMWsdMYAPJeELO/vndQHus9ArkqjUV6W7xc
5azvhht/2E8lH7ZyV124iZcV82UzCU0wdvKQ+UiNcStpei5BFE13Lr6roMcKzIqKsk2YKanK4vZ2
Yvx6WjzscS/eH6N5BaNvAJKYgu4B/lRGdEJVrlzBc0qSA1SGgjH5DelcvwT2rJrqXOmLBSYCQHFR
d0tLDRGw7+/2vK6vua6En7nCQXCFEa0jqYE6eJV+wJSYE7dGDKYY9TFjD2Jfcm2Z2jPbbCVjJ7L7
9QHowK5ti3DVPIbg5V1T/aZwd4flCskdfd61oAw0pGVSDPqZ3JyvgPuNTiMbs2NAfaGOA/4ds9s0
GV44z2QDimwYfth8vuh0AjnZIsGBJXmga+LnSF1EKrMpmITtpJgDu+1HIqE8H7DctzCssbh8ApdH
FO2NzPJ+5NwGfTnHCvQ9/B6Z+sggebTQHY3fzQdfcJR3OSIffR6YnvSW1/XgSUa2BVcK1eeTElhP
5ydhyF+gMlfS9qKUNAFvyeaaGI0PB+6gskCxq+93f16udDABcCbFYY76Cp6AgIKO+pa3vFDF6II3
bPVTDLvgQsGKGvv2pmNpAjN7lP+9q95ynI2PqXwL5jjaKIu05IUoh6j4QHLUodjZLcZgeQBQVgrz
QMRPRAvQ7h21f8j3pX5ow7kXGnr+nTm+y0hFTHSzqnxMKuj1Yf2r540CLf6zlQ1QXLM82hkEXRTt
abS/TUJ+CFQQU6WyxgqUD/SUzkLsmE7lSCbJcouX1S5Iw3sXIh8r+ysHEOLDxw3+S07wz2YWeoFY
YE0JN8wkhNCV+kXPD3B4iW5dEIN6UBWCpNe7ysLbLTZf7ShfeAQjto7ja9kAPS9aP2DC2vYQkFtw
Ez+GWrIquRDIGcbMkGKjpfVfH7vrYcoq7FqBUrZXBX6npwt2bR/7Yl6s66xP6aGnw0J3BrtLp4mu
xe6FVq+KtjXoaDZxz/5kSJ9ovuy8Zr+dPfftUn+LC1SbjZJPvbW+En7s3yZeKgDZllKWc8OgZuJM
BeIDaKUxfQf59NJAmmfIc9PrwlzQAs8ly82XeRFaHldKJKvCb9mhYANuUHa/M2iwRIDTjG+HRJ08
muILG3dl+ONe6rPlWnSblAi8lBQdR2ivnEYDqMafyysI0RlEinWoVEKqpplD7ZNFYKnK+oCPNHqM
M973YXqb9sHC0swwkA7VRJqHgjLvstQBKceWfnYMYq5fgYFB2FZ/wId1MlaoSVElD4vh4wXRL4O0
zFNLvCR86dbOwpC9ujBjmnRRMetUvDJB7xVTjaclOKNKoeDU+s7f8AQSX0PIC2Qh4gkJ4/1YJ5ig
inMN3kC6AbeRpbPkfN/Z/f57mKTDkDWmuvFMMEg7nXpC9NwZ1+M5+TCI1WfTKZnn6on3AiVnMjeg
JyoaNurS3md/k2HLKFZtwjE+grCExNJ9qwbNa7nzjK9YHN89wejo3qSNZ6S20XRL6wfbCcsANeHS
yW1yReCNE0MveSJF+MYam+5/tcRoPVGAttdxZjbCNFBZfp/GpCgfjfryZAA3dqi66GtN7fmD2jA1
d17IosHQOl+H8LbkPRFKtEtGDC50pz462V4YdFV1ZPE40gcoimU6KLBBVT3yrazzyLothMvT25G7
2VO49tdnXJ8oAqWqnLyCaQx8PwvT1OmJ44MhylsoSCT4KA9sC6EH3KZbGOn7QkWZVbkePjKWdgwJ
HThlLhdcBNqmKGM5l5bvITrtZSK/FpAApe9CSJs5MRCvmr7HxW14gawuXcpjeIHU/hdgSytLmv55
JSHgNGaHXelpgAUzE8q8asW0bB/Tpo3VUd4Exw6AuQJF7Siz4H2keiszF70AJc1HCobukVVXxZT9
Yt4yN4D1vQI71TvZC75iV9j2cWWGiq7KbtaopqF9l7qnp/6yzHkr+KZDujg+io424G5X5CSsx49m
fNwfp5fS8GsWsaoK08QUchwgT9M0N3aLsSQlUcfOl4VE3bKZZ7D1SaZYfDJ9Nx/4vB79cMwu41OT
KEFs6whtgg/W3SqG24toVs8wqL0dx5JdUlQD2hUdEKKAhcpltq6w50xPv7bb4XHp4idQraSQaKFE
U9TdpsTizQ7UbH29R1jK/p9gvqC82yHmdp+lIwcvhNUO90QCj3UnFWB7slLqMJt4Bc1MwmJuUtQ+
u07onHlCuQcgytK9AxjbLE2l/95bcWCmKcubIBlQPFzn6Z5f+CYibX7hxI9wCK6D8n8MYSm7EwOf
O/gZnCtuaLrc4K5DH3nT797YQ6rMy2SXOiFbfs9NtCp+oPsQ/se6BHgL5xFkHWjuay7VryB50BsE
+4zzR4xvZT2QhRJjsv3cdVSTCpRhV4Sexz0GIsETHZ70X0zQe1rjxMPd2VsKJ3DIA/pvQkgngA8v
bwZ5rIXyXpeGDNrP81w2+IMsOzmeRybBQ6p/h2NxS7/cNuW+XvTyDuSu9i3sPCFG8Ttw0MnTY20J
ss9z1r84PXHHPUf1Bjg7ZSf2fdBR2X/eTLNGXxV3JVwzlUPvNxYwmKXsaAbKptfGRch6ePuDCZk3
RVqUXbaBB9OSnq3JlPdrGhRchDZpnnjdyzMholx4bn80MNmS7Tws0SMgHyYMJv6yXFRrQfd6bzcT
N8LwhYkqf4l9+ypLhmXLKpF1qxQQRAyqNAycn2a9xWoVPBUi8nl3sHlIfhnAnZuLoWTreVuMq+Lx
AzrxkEmsAiUu9VoR8CfptDCDYgvJk6ZYC27V5oIpG+uBX5caTn616h93rG4hm37UbVTKEKUaPl9+
MYUqThRtf2QEHuWkk2dStH4YxgHSWeXwgZNqDWeTRgVY7jPnQuiAuZAURVw2VN8bJGiIKBFkdQF0
P+lSgk938ANIW5QlIAoNo2uLHqsOsOsjrvdrvW6m3KzNP0Vmuur4ilmKI/sMa4irMauiamQB06Mn
OT+eACvhHYjCztEA8jbVvplui4yuFYhu+xSsforkJ8+qDtVOdO8MmWWT9zERwqn3tTXpf8wQ+Gdg
sJGQKi0bQIDIUugKHfqAntc12CveiqESoXvDrBFbAudK+wtuV/ACnBZq3EOV6Re8MapLhcM/rllQ
gqhsCN5VXkG6twK8ati6hCusBtkbmpIXq1tpWXsr2pJeO6J0LN44SdPzBqUYMAozC6LG1w4nOo4i
ofN0k8YPaxdKaWLkhOkydynieLub5OMgm27qId1GXN0RBdYt9hA+UXWdD4O4EbDduJYH8+3x3r3d
XislAWTWXuWeJNqQNEOwMxGZ8je9LcosS/lfQKZFthC+bztsdGIYX4u4WNHJXkygH5hn78vvTYgW
MDTS8cy6qgbC9TWGna+wr+z2AiX9JBuTup6KkvqQbEAX0ooGurVlnZ3MZswzWLdGin4wJ4DbcgYt
JOWtaCFVrOF1HK+FOSGJpHzixDzZot9OX0YOC4Yxgp9R51OtqPPJWJ0zgXCmKWv+TXyWVHgeWpjD
LulfTLB2EsoAwyb3+KI6SnTY6X8s1l0Ggrx2dyn8VHkHdMAQBv8rzcOH3ZmOMb9jgLkAcPxrnKEi
fmv18Di3wcChPKE9cYe2qMNCwaG9khSbaiW+76SxhIcbA+eBpC3wsSjvStmeHn1chbum33cF5078
USVUAriw3qx/IMRutNjrU1wsEKAQsEE4gPri9qDsCMQJbXAgNdI/DFbwJPTlPBf9wQ4UJNT7+8P6
mFSTjNOgq/geG2g8GZ8V799cK7DZH1z+UvT2FeQqQZo79rIm/NhvAK39XgVRVtyGSc0n98jjYmlj
w8yfwvLmXK0JdDddcW3VLXsgs7uHyUhnouZ4kYIxq0kGVFsFc4MJWzEq6GfbPHAggxIB3CeEEI3o
cNAFunvUzpfyQHRAt86FNNjFeqZiOju18v/VXTbINQTGJuxy4WLLtzCJB7OlVmo9uuEvycO2Yw8Y
JticxyqOx8cG2dGGGA12EOHe2AfwCdXhqBmlWX7lxQS48hn3nogNIj2NgjMMa5Od2TGmzMdnqbGA
na1nUPC/M36i0DEEQkstaM6hnH8VMmLwK2aaVirJ8j2saDx3I1qxvrLkr18uJCNoCe23x9k/LfTC
5yUtx+eh5GLhndBpLW1tEugCXAgW7AQeuinP4qnVufF9wDfASDT005J/Z0MPSi9aXb06JUQyvGq7
Y83DTxT8mJJXyCFPNATc2NpZDWip1HMSVbQv9YG1fTKHOofAOZYUl3v77uGju96czoFdccry25XF
2G8/F9hBNrmMf0wBSo76cuuu0pOpZe3JENm3Y/42whKgnlsIriJ1JrQ3gwzVuSl3AQaeXoTWwKGd
9E7lsL18UHfbEVXoVeXG/u7Z1YyIN+u1Lah13uGGMSV4T9kaJIjwLba4IwJzARDafYg87hUQQ/bA
sLpbnw2rBhrgs35yFvjD2f5Q9P/Zq9uVRhzdbTio7tg8bFqMDVWibr2w9tnBSzQve+BkttOfTpes
UG8gP2mhM4RubpmmjHNcYQZvv5qDN3/0Vmb7F/qpOzoquNU3BTQalJuqF5OqjgmY4iDqk7hCLlCN
hxPejPVTo8VZoZ+jKI+/3TIduGIdr943bcFzEL+QBORSA6FwCozsbnRGEaC/wMdBzPM101buV5BF
hmbeZ//kNGn1E9ldLzzGvFvWBRAmbalFAZ0Fjdy/TQ9ZMd2RgbW1OCchEp7Ayu6bVA40fMF7WvED
5XEKVNAiLjFwnjzJgyL+vOPYrs+frKVnfo3aWjIIFj3YI17dLG/uMZb0dcEiXDSxnpGxbBr+TKpH
0UfXwlFm8Ox2jq3v7E0F15hjJFxEUcrvL1guxE4+ju9m8G6VEA34L2fZOEwUdz/OCsRmJDHVb1Le
t9KHqxsota3nuwrzLDRKDEXtFPkzcSL4boGmsj0B8rMjk7WqCHWvTzaZp2nX8ekLQxb+12jinp0Q
xQ8KWmKA+0c3cNr0m86KY3iowHSTA/3nKTEYHGVKOhI/aDeREiW9AGTPcNDsdky/fsuJDhv66ySk
ErezkDxFgPHjV1cK917SgrV1L2tvB2HKBJUqiRhCeCT7aCbPWSC3arIB0dLQir+wgJbUqJv6JZIC
F8Ov191knThKkR2kaY4h3Os0qknNQ1iFCukz7td5bwvhVuWF0MgPVPprldoa6COaQBk5BX5AlbTz
TplLsthFtwzTaZETSX5yReCFCDXppJhVmoB9Z+KdUz42ny5/84y21N4i7tNFYUMC8xav+UUMNrqX
TAkdsSUQXIoIbz1xSdCXbyNZLA6p99f+Njs6KAQFot2QDF3bV4RtTMWmxPx7vkl+1/izOSINIGvW
ln2hZDwYOH7Gx8dhHcuFNrNG9cHwo8NYXQ++XJcRakzdYfE+7aAROpJzykAccEHkQb94hP7dPVTn
Zzqz+7I+6CmlB8aAiWxTU4ev16sTRr/JDr/JvV+gXwSlQJv0GL4mFRT3xQyQ4Q1IQEA3eny2PMWy
m5VgLQLh0R2AhYUzwxuw0XgtNi6d9quBc8EDI3AYitE5qVfOYWClfyIqiBE+MEkbv2uTImDOLKWz
BAfqMrv8cJ3w64OIhwwb4vi8AlFTfUXqBh0HVqbnyJj/7Oop+iirShYOBouU8nI3c1qk13D7a5Oz
Vy4cWk2C2bS2nx2GxozdnEewyArUTHjS9xrzy/95z6nm/3oHUVe9Z+40FyyLrclFBIU4WJK3xfHO
Fhtj+lXzwX1X7yccusVZAKK3e5LCVQJUyUCS6936T1v1KtmTq8xGw6CJ8Zgq+ZYD3h7O2h/w7jRH
j/E3tTbvhb2dr0tgsaDXN+N81cGVk4Pn+Ue43dCZYVqesvynKG00zCibqzXlBMuVKJtVjINafyQ0
7BLQjaARCFs6HFHD/dBOYOvIQxh6x5OUNqHXOsSHI/aeBHntyuBP0ZrUsNTzll+zF0bZjD7Zau3l
apBB9XtntTBwOMJF0cTxoOwTD8CAtO4neynYbsWzyvumcBaRc5ozwqt8faX2fcy45QrQIZGmBUOx
pyKJIqZULbruCgRfMtGgQPBPUaXWRgzQOlTpxWJLYpD0L7V9k4jamO8KI8RjF1RxICZUJkrYhG0W
O5u3+tvXML5d1wFpUO2ig+FXdhQZ/cMAXCv7sX4xoJBhXDU2/g/QowlKZ80J9/8WVhIgg3c8JG/S
3IopMaMzrx7ATA8/gUfJu99oVqH5x/yRgZoL/89/hddfdmedgVFgkPKdlgdX6opSNc+PjX3PX+OT
RKFPrOlGPWoX5orXdLm5+0zZDuzUf4m+Q8wp4+Rjbo2Ms0o/SYG8rFsrf4zJVZobVjYAZwo+LLxe
uwVwrG+A/1KmqbbBINezMGfVBZKy9xabl2IkyyLruYUVDl2kPSYCZI52+22P8ZikjmiWcIOzV0GL
DpzlLKmtQZk2M25gDaWCARJyriNu4fpN9cY9o9nn+7L+F87w626nCDoYRDP7CL/YVhwjD0CQn3V1
XsjhjSt1ushxM9vNmjWde7HaJFVsSnO2keDgTgUqHqQ77qPxkyo//MZl8AiuAl1PujdyMZUC4A4Y
TVUH+a1Mpn4gAdLfrq43a/S918XQ+tFyBB4YHCxZmzMbZfBZKfKry3LsAwfPIzLA1xAeSMrp5Mdk
/0I4hDQKY7ZIoeqeEEmmq3vZzSLUk/y4rOtJ9UFY36swQEX+dpazbUZEXdmrpHj5iLTbavhrSN+k
rgl6S2SiTb405udBmJ7QKerYIaq8JI2tsazcMZhnPMSkWBOC9TH2Zrl2atznEMMoVuAMqlXLvYvk
79p0PkziEf+Dzwriu5nuf3oTLIIfCpPImVOj2ouib8xYIzxO96BBhsWtPrfT6IxFdss0kgKQEde1
G52aDeKLtyPdj8WsispocPl00IKn3uun+y5ysMsDrzEjS0GwSHCdLS9bAVfPEThNcW58gWwMBqR4
2BrnUPlTGdIuDVBZ2GNA4HK/h2DApk5cPkH4puc3BM4VgArXwlT2rBWXSe6VSrXmx8SnaRckiz1H
720BH+/C80lqEnFQYiQ/Prna+XwyogTNBMIHvIn8k3kGXqGWLelBdowZ/P9TZFqxRMc3sMbNVkS9
wm0lOluEl+JTBMu2VvdePoych3DIwIfLmaygVKsXTh3C06XqP2iU+ul/KajgRLZRXUqZ2C0hSEXN
Qc6MgpF69C2aSjRwlA4iLExQNjPnVkkKDKV1tUCIdTIHmqA/UMetImkdCvIM8igocWWI3bWSJeww
X95h1Gs/cnBgPNwVcqgoNmT56S9MGravqtkA1GwC/M9vJyeD0Mt+f5zIQFQPMEkMBm7AQFg9Xj/B
x+BiATkrSCWPtEx/ttYBvVeL0Hp5ytEuZPe5LGg8POdSdhcXQPZVymEHqUgAOITLJ3K0iVPwu9kK
OK/6BB+RI6ZOiuNocZGiFHaxKmb+gBA8a/1/qs8pWwIyuTKCYRnDP2wTJzZ91Jgf4V5BPS9XTmIB
AkA0dOzDuCv7AFT6QzNK6za4NWRNw2qlZr0BLmoF/ZcVMvFEMkpsZnu6Yp3qIw4uB8+bwAzZilGZ
exYuBY7W25QdoLvcBFRNUPeKE8EF6fuqhp1qr/kl1TwjT+CjiWOwQM2b54NDZSeEiYvelLIRfRUh
Lg/qtqs7k9lxbk/eBlDc6egw6jPAT24sHLy//pVjMFyrHjC7BNZksY++Yg6OYSjKLo34XzeGe0ea
BhgxwI1bfpasHWftJQE3rK659vw1qQVPT87hw+1sHM5EqjKTD1cTrANDACOZYIJZmhGN99HS1wi3
5GNGfSYSMHY/VgdAni5MTETm4HMvMIBkKkoywDpQOOnSL03fW77iK8F60/U8+s0tobAUTJve8tNL
WtMkDCaolbCqMg207+4oWrvPmtDLWba8QdEcZSrJQl4bug5z2W85I2xzVY2JnB8DA5YpwrqIs/LQ
/40/O0YcGCwxMm03qKr2lNVKk3lljyEguen2ja9qKN6+STwPbqDjpOdyCxgUa8GudgMg5YabeKMt
0pBDWCGaJMoZGznMl2v7Ya9CgTefNdCjletzb4yDkdq+KB0skNYacyGGLiyia/DivwGzq57++AZX
KJpuNGavA5+rBcnNJmTu6wWqVv8LJ6o+DHznF1+cpwaE8+iYXQLMCha/4vnUYD1EhfTKf/EJJL2h
lyDct88jystF0xtJQEzAB/i8IT3ERea5Mf1AL5gJGgK1V+O1b2xQkx2TIM4WwPxf6MH+N0sLM6qt
XZAyM2QMEHYwiM5ybC6Sc7iw6dq8mgJC655WfiNPcjTjALJi6vydhnoFj6IwZhDhp7QO80NLiTP/
2U8WTth92h5HLjcEn94cvofgYQO9+OCe44mc8zcNZYk/+sJO2Fgo5CdxqPjPJYUJ3ku/qQFWYyLk
YhDMJ4lXqiHPgTHY6ZtIBYDBUrrtehmbHILClF8Dt/FBVa0M3IJmdAQ1wzL8g5+3g0LglpmZbl7x
o90VLttBtK0cKf7TK5mOPDb1R8amaA7az3C+eVzJY/mtgu6wn7fvaDn6DmHgfVQkuzYmUOY07Fxr
+S6x1c4qK2udbFz+rpAHLqk9scOD+H6LUSLftBdX6V7vzZ9moT58qrWWJWBFou+MdaK3pqsW6GOb
WJq1bElnxzvBvXNM7TG8aCY8Qgmo36HVooHb0vtFIIN/fDd09XprC7lAJDYp6iOTfLlytY8O4TNW
oCR+kGoWcVhMsYSHaCi5biAa9TBfZWhkf1VohWfFQ2v5RAHUGuMRAOIE3VpDadWYwEHWOPWVpqSn
N0IDjyQYPFFEqmwGJHCk9NRdEDuq0Tix95ctDUjIJ633wIw5Oylyh81855CNd2Y8bYArYWni3trX
jOesVU9vjSd+PYHB5AqNerv5n0NE9E2mFN2BfcFe0uL4dMQys7+A2pPAbRmCqMPlSvmDHHx17zCt
4wllOmG6sCBWfvomIj6ahN50SdbgcEq6/CCIrBVNnWIRTRGKLGBT7uEheMkkudJGRNyT9SDYQGoD
byRt2JShd1icPTtbX/pUUiGpkLeip34szi1UBFIwceapJcuL6FM4yPpl4du4ej6XkClbb+0BbHzA
RbWJaGZJBHpZf0Oc+W7dfAz8sYxG83NZIsPi1jKNyG4ZR+KJuzE6BsCuVOHn/7hIHZhOADhZodlH
zhHwD6E9ghY5bduoHSxxx80r4jAUjxz5bi6F2fikrs7fj/LhP4VdVF3u6naDsgzK5+4aUEH/CXiy
Vsnt6Q+JS6wFQs+ZOszlZO9UslW9AMfoTmeDxFjDub21J03sMJVnUVnU5qzDSBO0WIwTtPLqaPon
+pxDEKDV5xYDJO5Bttve9w1WslMJWwRJkcqjW+JQ0DSSYkODnbE+BCw6Fi4yzaTBcL52eoxROVm2
pRMazIvrVwCmmgC5aUBiD7AihG+23GAC/YNJtdmBAYDgOu3QQwv6uRgLvb32tgfbtLlu4d+VbeJd
OuCe9qOOzxvENpnDUfdTAZNV8cGRLqWa2G6j07SubOQfyPHl3qYCslyz5QmhQXxUrnYwctwmFSAY
eBh05I2HNQpFCDXo3ets0tNcO3Zvdc0JlYXVyxlCr8cVnCcN2A9Dlt18Wr3hESkFJgwOxOy8feeM
IGXdKVdqaZj0FdSIora/cNa/oNJSmnGw8xyMStAvn01h/snxvQIEWNRKMuP7khPuHKOZNnn4X7N5
3zQFcO18SLgSAIToqp8Q04Of7YdA+sSGhCkMlZafUJadQrmxIs5fMDexgSp8dSwrjfNqmAeUoeLd
Iiy4Fq0Bl9BTjTTPbClyt40syx6497MjhrIOaUjRCheqGaKTQ0js5D85AHTpyAxBDDx1ceRHuaV9
i2vQtA3Kt2Rtp/GbmGWG6DpwnMIj/v/PY9JfQn6LscomwvPMb1mZOg2JPjJ+Mu1z/ZuO+qjMnOtm
wFZljy1Bw35OF3fuS1OO7NIjyVbL7YFmKuCafTtr/OQP9VfffIV+OvTysrMVur9g70L+4t9mS+bq
bEwUkEuGFV1RnBtMR4BU6GvSP5Nsveb2h5xIDvFZ1B21UAducditaAszJp9Vf9fseNp8ox+6NW4e
/qULbtR/wSW46kOGpL1ZP3KNLl+Ok1cccFVXyFbXSv7Ttlvn+eyJ7cgKVIUvdDzzQZCd9uvYiHwi
PK85PI5miF97AC+6yHKMJsXo0VNi3nehRr5NqHsUlEVbw35MjHq8ok8V7YI1hq/X7Jb2AcufSL7I
u++wNRDgWJ3JcdnuZpSv1O/4quZpLNrjNF12wmqSI71jCf6M+5TVFPW/yse+L7MaiBJ2D6w+S2Kk
n92V1Gk8XHP4fIoLzlbkUozKRpj65LQmlj3qg+rrzAkQ/flu7zIU1N5nXN1jGqQBjWpMFdwosO2Y
stP31l3sjM2B/mDipf16PboLlDOZutKyVHvzp2PlsqqHsbT9MT8t5YO8fCw8hEFFsMGdncnr90m+
/q6MJ9XITis/0b4//1nSejiuLx5Nndfkw2v6LJL1tvusCDM8ad5iNRFleqAaYu8OCJtiKP4Ic5Nr
F4U8AEijs8Ha5o339hlb+hsJnKMdfTTUE1zBU0KBQeR0RcDxeMfijgEIhnnxXesahHTSqwIQMb0d
YNcp8Sa3meX5bIjHvS/x2PpJw6/Wb5AyFQe3ZC2iMvG51QwsEKOii2XPEhMqNmfMJq01XaUbEfo7
jNhrq4d9KAjRduwBon7KiA2ZLHojT0eHMv5OfW6QiEHR55rNU7bvUDtBZBZ/wQt1QKoIc1d1r2fB
/ej4VueYiY7RaMjM/o+zedDbIJl+Q3pPz1paceoZU7u1d5vrvrUtzbBsXrBg4WgwMKs9W/3ukJbS
FHXhs/Lu0e88qA/qxBLzorPm31WGmQm2n0Y5pCYPkPoi8j+tcA9jW2oEHzHts4Xoc83WuBKmie8x
tUymXfdPfjioOBU/Ei9bjWNC3BzvsrelZYsDam56pDTEGK6eyL8rbISFNa/6o5d7qaS2c+VsXtAz
pmGizI1vST6ojWvRQAKr1Metzq5tmmBlSiSOfbnOV+4XlGd1bU0AGA9Pvix6Jhygp/tWUb+mofdN
derR+o0RmVrBkJfrFRFdS0QxsJA78pCF7fWvZP0MUGoNqAlgSXwYETqAWP4o0hrZcNK3Q1sYzBxg
NLS2f0OMPZGfBb7o/cGv1XwMspEQG9k1rW4fxHeOvSIFlNGAzqCn+NpWgkBa8KJ2PwXSEFERWTem
FX/J/dvC0luHei0a2zarOu3qit5BHIKYSC+67UoCwpXUVo3R4NoSD2+/Tbs2S1SgXy3N9s0sZmkM
mx84x0S7XuqWpB59e3WpiDUjP7gdMu7CL1rcCwDQuoKi4j8eD6PmY3RxJQXja8xv3B7xa3QvEgEg
Cc3MX7zZW0GmPfkED86ySXLoiXdkEi2p8NpWVl+6Ljau02cYAZTq0UZyLtpMC0p1X4nBp5dwBpha
G3/q/cJpgjetElTIZpUSqYxTtGQd1SezyDFOgNyG8d/ATdEzqjnFfsb075dHyLd+hxUffi8RZU0G
9w80ve/mlUnWGz8+EzRMVSo8jOYJAbXZ7A1gWVBwKDsChv4CJPLjF5HeH0+28uIdwE/fwyeX/5Yu
3XRRIiNcVVyWBcz+sm/CUS4gclADNo706mBx7Dnd8wfKMsAGjR8hh0pcnBQ6fwn1js/B7HyTtrNp
wTTqxVc3rOieHpvMqBZUmx4darrpSgzDFKZCyL78pMFHeuqbgRrL/i3+h9xlNGr3b7SUbO3iLrZQ
lwJlKNmfO+nKVYhZwdTCCyCI0Xy2SRodDpb0KDibChZWul8H2u/2qQWx/QdEe5O3xUzgr0hlQpCV
mOUOs1/HDkPsbL+VCTYmZnE01ZWQ+q7BSL3bRTBel2Un0UtdEcgTnH7OEZRtXc8A38pTZIH5jRzF
3UUbrVK8v5v0IVWORyqYmEi5Z9nll8L58G2EoWnuUzX8D6yYVWaNMjGEn4jvi836ppgr76u0mJOj
lqPU2kjCYEJGa01pGb8i6t0zOhGKbGWOxvbExC2Zj9U33cKmRR/JQH9Vkj/kbxTWzPQ80dfZ1R+H
+CEid7MIWdRp+K71SFugV30Xx0zdpq06xn0/simsMV00uzpFAXb5orqWnyCpZL7vO8xnK6txmK+1
brQ4BudAspLWxbTmrJOwR0Xj14RNSiq+rmIZF6+AYGyugOoQBMYArx1U+qn9sxjf/CCpybqjy3kj
m8dbt5/SZY2q2j2p1a1UaPGB2LhH6WvLzLDLaSU1pC+2zwbJnDJbUMC34BcA/b8PPfSV1nqAt1Kg
T5xPkyLWYLy54rQMHm0aUnywQ5klLlNvScq35zEc/vpoQ7fOBPU/xpzAggMSAYhjjWQq8Qw5ZIL0
QD4HHGP5nREJlkm0ee2pKah6PzPoib7UHN2QuwysFjt4m7f84HPdsyG1iuCWXtD6QA5HMq/pavAa
pJ0Kr5YfFQjrHCN1knpxzTwhD/65kxek/RQg7hgcexEWAtKLKIBahMqGjEpfoHzV/1fGJf+/gmSc
Emn46hV9LpZMSElOHtQaVHk/NO079JYEzzfbfTSCmaE9YzpXkEENzd7RhWbqPmVrOCKBkaJIE2Ju
S9ncJa70Z3anD+xWkMzS9uZ9kMR+YwTYCgKaYIk26NgJls8CeKesoXiXl2tjfmR+VAs/DuQ0mMXy
cPJVHpaOxclf4tiW05R/3Zy38z66noz1cbO9Ht18ZEt1ewZVNJC9nXsjjdQa8OXQQ2eKwwsXlQpa
FPwTHGrd7OOBeDlzPNzFD2AlPdmF+ouiq1KudPo5NhOA4WvTwYEvWLzHAL52RoSRalf5WYDjCTt4
sBJJJCq138J4vspARc4Yk+uAOLMMXFlgbtvGiQqfkUuz1Ch5IATQl0Qcoh9m2zjdI0Oj4ldzvrEk
1PD+hTXNmoMY4LJCIPU0wyCIQV8keNfD2xDdfhxtcqIX9O6N9GrFEUKaOO/AADd7VkhXZocstf5N
F3+UrA1Qt6tQL9D0lBzDWFvFeAV1bK1XUu1lQ9xMVJwigObTnspb6YH6Y+4YdfOCKsduQI7d9HUR
mM0VclpIHW5DxehZHTw978WgOxJPr9dYWQHgZOaS5GdcvTO3v//p64Rqhl+oNoD4JCIFHNAnhy4z
n4toCylk108maSFAQ5hEY+kvbMRNe0ASO+7vTXTi7Y6ENsYxZZDGnCJM3iCg/qXs9DZo7M3bEGlN
+g1HqFZJdIK2v4d/gVjQITdEx8s7dGoadT178nA6uhnOka996sknsq0mFesSl9QKagKbY/3QQ9+A
+NaD+9yVAbNkNTNrnTrMYUdA/Bj/PaaAH0wcSseUP545MeJxZ6YJNcgLMsW8wbsvpsmB/9Tp6VeF
wIykKuCyaWUupSZyuGz66NTV3dirU91FxSas6E2Ol0LToMsmPppV7LfmBvZW620l4G+Bx95cWXhi
bcdU72cggxr58tfXw+oZMVREh16/2nXGPqpVbJ5CAK+HzrULLcqQpdLAZX2YSOlIMHRgO8yN4xGB
BxLZiagfqEp3AzLPzKEigxb++C7AS+PZDCyvfuM2+pQ1t8bMZstjIFI+aLzKVQpDCYvqEc0hauch
i/zcaqOMJYmtnpfM847x0vBpNDVpXwyXtmTzscBXfikb7yaKV4V1h245n4PAR4nAKYee/e5Ojm7S
kyD3aM0QLO3ujaMgEj7rxmMBqUAefwXoH3K3m/MEuolAbUcjKoDWjz6vGn/PqDeNv0NPkssn9qNA
HxF96ZD37hDs85YzEedIB4ZEhwmtuj5n3b7SRmD4WBjsfwfwfdeJE3UB9xPo6Rrb9mEGepwpccQL
4Dp4VkALDl8ApzfTQP7kRZVHl4JEqWig1zEICd3ew6QtDX/3um54PjGDffoSmt+y+/IycQs2jgl1
hmzNhaFK1QOqKEmYkZIVpkTvDNWqHEESR/6LTSlqcY+Rk7TR304S6pV/pOpLe0o0AiHUJ/6LSyfF
POoUc37HJl60Q0/lZTKNyDPzpFeKC1YAgjoXzMDjnWQF/CiHUM6pHnCaOq9rXaj4ph7kQwUkfIiZ
3tJg+XnSQuOGnhLSlLJMmCdY6WeeTqzRQgGRFGgfnVOfEM8MEtfTrZ9OsPCex2e9cqMYwzAqvx3B
SjDgdP3tKDUchVuIVomkbAVJ+exz3LFIc8jdTwQhcXi6kz+U0vcZUhoEVNQmjf66PibvRplOXVfT
xKD2DLu9SXcgyNgwvY4a/TJlNSiVWqj1SBURkbUBMrvRSVUH17zqfWOcLg1Lnrf7QFns1kzdKpzy
ORAl76DP3UUMH+Eu8BY2gt9L7ImrDdcxDttrTkAE7cG+54qYZy7DRNVQPHeT6p6zXmWmfeZ98+qg
9opTx9Zi/yn2clGgKIFycR7/Dx535s/Cp2JfiY4gAxtsyt7nvGwaKv5xfY/fPYCfDM+htAPRxlUP
kpyWdQM/E3fpEUhhOzB8U9hvPdGq4zaUULT43dJC4km03grMyWVNE3i3MVy53s50RzcoJXWoY9K7
shTY5CMn0MU8YQ6VsvVljMQ7LtGhWumvaICwOnBfMzbjMxyqh1WR0/1j4EjAANSsZ1fEa+6yINdI
csLZ34SJVVf80HturiPIVJK8GL4pAtnhPo/FKAiBRUwFK+myHAQre4Pj+00CftYAi8S6DJO+A/YS
rJ1P3Na0EN6YAikI6BLl1JfLqbd5X0QE9NAJHN8w99rl5vLkuIqWRbpRjULUlMLndSggBkbVbUzf
H4MUUv3UhpFfIa52iHRDM8O4MXCFkxT0beekgLYqFmGbLL7W98r//4c428DRuOiOBw9/xZc73umt
8PUYFIdrFpLMt3pXRbgcd3AF3u5UKCtnhXfCkypzf4x+U1ToLLlN69GxOudT+VBmDhuC52NY87SR
4ji9BWOJLoYQYy8stTS6JcoviWa3ycXuEwuGYDlJ6+c4aFNceu302CQCuT12g4l4JNl6LyR+72Vh
VlHoxqwUmFSsFvLwpudl7G+bL5Z3WkvZaAvP9tzPPAHxGw7kgrbYAtDVdGU002TNrfNk7TmMOBkX
8d4gwgLgvJI6tFrBlJPPNs5x9V30O9zBHh+MY1YOO7KqFFTKCmdUjw176ZzvbRoiOPH4IituWFHG
CulNlgvJskpMXvZur34Jq7EV/j/Wqb8Vw0/Q0AivYUbZC/0dvuKXY2rusiChxCbO3OpGjZLYOMxu
0NCOhNxNAsLGIvLHXuHyBqoHK28fMTYBJdqU16iZEahwgwHWx6q6+yeHgm//CyeK/r790K38SBBh
YPEMOYJSvd4lve2iKdGSRYm/L6o1Kz0/qulMq7WKInIx72l+uhXduiOcLC4FmzusseU2+mBY14fz
aoASCDwJ5tXu0SN+YIYRWz3rJOp1Nu5GKAGPs/vMn1TlWCUxGgQf5/1tVaRsEj1D+2daAeDu7fnY
BmGZ1QDk4Io2d6Lj+umCBD1aELqCwDnkkBK+ge4f9rXAXOZ3m3ZNFCdpFtHAvwAdue92SOLjZLlw
TVgPRA6RLEBu+awHuvTKU6R2Zota5oPcjdZhs/ouud5bgtieYKZd+57kk+4qT9RhVj+9LLsmFU6S
3bnhZaGgv5R0K6nanLPWjEPjDOF8GQmqnOKBUpcwBPaFMDEIfuAZqOCxvv1c5H9g18+iH+cf7cHs
lLgIC8hs7rEbUpOYSmgiQYocVy0ynql3zHRwqLUWPmV8q8THpoxyrLF+FEo4OjM3tOh/823/xLGA
3i1xY2+bvFNnHOL+51nUF/c3mDh1UNTrCfAJJ+20MNjNxa6K1w62qE4R9rk3/2udB5iR8Pi3g8g8
8MwKsv/a9coVCLFXjRKJF4T0CZq33bOBTFHQmYEhruBF8ysic1yf/KJlJhozeb/h6Wfpy4T7h1Xi
9Vx34eLwza5KIlsu8f9Kcm9G3Q6VoFkUodJlkKCJ5kTC0rGA/6jW94XSw+OUHtu7gdnbbIHywGnl
45Je0l0AzhxrrKPWsfVHSuEi6qBZoXYO6vB2c+J2Kj9p+bWMsIb2xyEVGWSrydT7525kDir4HYmH
iP9QS5zgMbLc8NvuU36YOmyfzEBWzdXWPj5evo6HMdqpl189d4PqMpKPc1ANHqF3VWo9rG1TuIkJ
Q5MZVE+u/fz2wd352w5TjZ7BD+5aND40YCPpHx1qhDChOUQfX3A6bRoeX0GSVyh3r4++Q9q+EdVq
+G/sRZa9cIlTeOCC+80HV3B/kj15c2ycVWnfgQqFrx1uFf4xrRgpg2m3r7el4AP6LnRn53OxB+WR
CWw7x4RMy39tPkP0ZnLoa8khzmOGkqHmYKiUOeLQQSpxJf5sy2ofigcvwiXq/MVUiTDJvlbZfnBK
Q3S1mVZxFve3HzC2J5tOAQ9uX0At40f7WIjmP1buRatYvTZCBnAZzmvruLH0FvgRnxRfmguwzs6F
QmSomq1vWngx2dzUfbyq4y7O3pwDI0FPLaH73cCyzPdsrgnkE/JOmYAOMsV0NfXO832rq9IyHpR+
ix03FJRxrVKNYrw66LpSchyEJhcgaYX2dnDla0vsrMrcebtZMHNN9scXJWM42s22RduJVbq5Ko86
GqMP4yqX6921LA1epErE0UzhXVM7BV3wP6LqLoyh6BEH0fewmtx8uqrq3JTTrEinQy/X/omSJ/8o
+44oEZ/vrmHLRG4bqmVY1Qkf6F65SCLzh4xapFgOP5Vbv2VUIVPpbOOhdVZpH02gA0FJxdbJUYB2
vtmwfrPA/rgcuN5G+OMj1SM/54JisPkMz2TmgXhYsmtzxeYWl1itqACLo1SmhqRFmLOXwlfQp/Hb
3duCmudsoCtS3hLeKmnzJmi1Rv/OiXL8jjVHKjoqGMaY0ETcVn/1seMQkwzRctHklgWfboIEbtba
2CNTvSHB8qAxcsio9cm+BEgutnLWiy8pFSlt+dk201i6IFegV+c+9T46iDhdBI2Amm+toVHcFsuE
w3ojIrYGCyvFmPpSuHhHH/F5zTVy0LIkliKFaLK9oXbIlatAZY4kuX9y1q9XtqGZoom7NjXxR/Fo
WZd3Oicp0/9Gfz0ididghZFH/vBOLMzU+LC3W6MlvNKKVUPYrYb+xx0v1l4xW+8IbNOLFkdkhAJX
/uettY/kbrACb6Bj5pqSALOdjqg3ytsShPkhXcUGHFVRe0ooEqNOSiVHrKFUwnfpSTZzRm/I77+Q
teYFj/6g43Ir/JCJWZcAsqSZGX1C1aO4a2rd+LAIpRIlVv+vdN/rwAJpFWdvsVIJTJnDD4LfszJD
8lfkm6/o1f41dtrGmKqHapLQRvPyql3o/GaqhTAquvykGA6+2wcyJfXzsnDd3SzO5DYarGWKXRBn
dtt2FNCBv0OV2wiMUjVWuYRZeW53tlT4M+IiITgtGT0PVs6wsiBh9DDY7gqqaRDt/T8Q/nxxtyoa
0MDsA/SYM7WPp1JQY5d0O8+WRnDodI126RHVJG+/jhsjP66XKchIlQfn+C3IFKn3SUSbygvkwmfc
qoez/k1kQRJTpkXihRSCwxxnr+OQUlkEFr83Dvp0ocxiHa1yLwCYNXiRvd7V8HzSMh3fXXD1V0O3
/xjXC66Wwcna7exSy+FDJtpwFqeosk9zz68VIgG1pUGt2lCdcIm+71ig5lcI3vreP1/eki/VVwfA
vO4/RhFo9hFAg6pc1kgr2GwqEaaGlDtSmhHXmhk8TsEQyn6ZbZXCwvazRalrHofnxnR0KzEUsArU
WpilSVctDxGePYb2qn7yKQ63tP5R8MXB2+xR9Jog78nL3AfGb6/+Qx8ZVLhNPrZnLGPUBE7dYcgE
jsx9GqA9wFa5e8Eujo6dLuf3CudvkyCGd2A9+PVp+AEZ/KlVd9OgQZYf2OeFpfTXBtxJgMmtqQJN
+IxrLwRJMSb2mmw3gQG8fZTczi/8IWBtzKB7uc6xBza1/ytCgD1ehOqhIDRF8R145HbnvMSEGvm3
uhLNdVfl0HIQirko31Rl24KNiRUmkYYcdpdOFjnkCDZJaiT9Jzsz9MW5xZmfK/qgUKwJV/0MQsaY
StjEy/lV5YLFgJndwcmQ5e+TdwGBH6+5YSRwsFZrnoeY6lPw7+ZMeFQUj+9niKX5l6aArs83hky1
eiezvhfCZIZUzoaZnFH//zSRUJ9iS2uLsIMoWGjYuHiQu7GdzwwFYdgrsfVoaaWkYzg8V+IqHv/U
BK5QOEg12/pouN/9GkTdcaxJqAcObovQpevyvY58eClO4KaOy4ki9KLMcRZcx7UbRjP1W6LYGLs5
PHBAsk5IagjAQVi+6ESvJHRoyu26x7Ga44y+YgqAIfTfSD8e26TXp9mrOY3pnyv8MO6EpT5zh0yf
OygtDak/6ZtXEuInNh4X2V+iLYgBJb07qFlWa9tFLQ09Q2bZd+FsN8XmOrVdQfwT9ityZUPk9DJI
LzmcRFN2xRzb7brUogYjAKv9T18itXMvszk68A6nQMSsq3wEKAsxWLdQGcOKIZHUZCQ36ClnH1Sk
0khkWvuIvMTQq0Pl9kXgRNO9/7KsrptjUkMauJISrMS39ZbcuFqMe1HbFUFZ4Ag2Ij650dBc1qV8
gg09cC00E/EUg9krqSp/MKprPLsvo3wEpEb5XOKicwWxYzO5HbUrivDrnujrNt92waTgBeP3AmVi
9yFNBAy43Plzf1oJXHs4nLdWvho1KY0YQ23N8WpK2+rqvBX94tdiTnRhpVOF1JUbHxzIF36KJ0ZX
J0gnOoGoR7LdOOEfoDjLeyclB6W/BjEId7gh5TMWZPAHEDD5DoUPuGS+uVru3NS0kYYfPyDg1nGo
HPIF8z64/FHKEfHIoIjzR1PvDuksf+OZAUYPZ9oFbYzBMxiX0rId84RqJyFibYWeqqqZ8vz8p4Sc
XxoQhIpHDW8PEPDAxRMgdjXbEvu0ICYqeqnM5kv715N/V70QfiuEyPr6DYZ5tccqN5YVze8WGNT2
jNS8nhbUMnd6lDEB25NCzBNdWvP9YF0rf1LLmecEevBQ8zRvTCCl/vlaxDXQXhLB/HeWrXnemhOw
+4ixPGK27PsI9+bsvTkEmP7sGXerSaidyETTVvWzo8GLqA3Xc2qbQDDgIUb8/fvJpJHc11UTJ6ji
zgl6kCRbD7qxntbiH1B66rSGrpo+TwbRCpUz4V84kuRuzrCWAeCYGwDhFor9JSQYgtJhvWvgS64R
v29SyHkTj0wvj0OTsz5SlkHiue/AYZySG0YPkRSlikNQLM1/0OOtfRbQvFuc+IEG2XCI+c86C9T1
2vY73zX8oka7zIejgaoDoYjkYp8BGmF6vaLzY8dwfejactBFUrh2KTXBF79yaYKhM5iZK7cglsZS
6c7wzDNUhs7E3Ne35BReNHsSQiQ2VTpqGBtPwDcSVhN+yk7ztigUMvsgK+AWAqvoK2O4f/1qvv17
OE6UYwPj/L6M/AcoRXqm2AxaG6dXDCXQ8NCYNjF3lBTSvWsNy6LukvLGw60Va2/zJ+EI1lxjdDzG
HhfkcQCcA4vunMI8tU2usqwTIRm7N/yCtAvDUXHr6wRJI8pYbMvqvlYcJxKQ6WlOqdfVia0HMF8H
DMKqZjHpiSAIeWzaFhjpMylMfAj2VfJKhheT2Z6dpu3OkodHdWXeiGVtO6oslxq9d73082jHHttm
uBl+/wPya7X3/57yehAttIB1kiFPelMaHQSK4vA0mqEZ0cE2Ai2byoFgdGFF1pXhiK+ITn6g+fvc
OCaCz/GGcGHQ1PxEiYg2z97BVsvCQboQtrEZDI8mLQodLxstHtUio0Cosm/4XiSM22Uo8bTWMyCz
c59DVWLdzK3nNN5jTh/8ktsHEar7qXMqfo6uVHd6z9uDizuIotOfm87x8u6Ygu/ceaAvxbK98/r+
2Byf+5ET7gDh0RVgEZW+W30GA53P4DNPlWImijDtkoynMh8hJ5JqIWVJk/xVNCugHtdbDfRY7nPD
LejEVKyKEYVR1/R+GIxDQ6O6F4+QpBrBURXfexjOs4jwJCJP/k1j7vQcBYqg4r0biV6duO3wphC5
JKEM0mPn5ZnfY3hDDGbjRnV/VG07xXQEyIz497tKFCX5m9NXBB/PN1My3/yY/tHjHJ6x37C1YDvB
Ksh4bOnR2dFQ+EWbKp/vtwOeAd0wNwB8ewTkQ6iMBroFgA3Ri13vf9o6jVAZxMJI7XVrsNwzbVY0
/5taruN/sAbHV47tKBZKPspQ/0ji9Rk3RzxP1egxIj0z0ECD2zTq5fZ3zXzSpBQ2rxSHZnmvF2UF
WdRjj/x7yrjpnfD7qih0XGUsBgLhQWqKuFHC26whrLH3MX7iBUmeEHnP16jm2GlSJtBLRcN82Tn4
CAETWbt2xyjDyYaAd8K+1NF6aaKRXSfIg7SUmtEfnNAWyVrlpDIZu5MJB/EMOS9LSEyhidbye1gE
BNDp95VnDa1xcKmQnyE9SEImagQE1YKQ27eGDnw5Xnoahkq/PL93LMVvtf66y+x6J8OsHparpzqh
HhXtGlydRV1H5Id4EAiLsiTAHR1OdP2To0d1XArbdsxoCaXLFWZfnZBwuAbiNneA3aUCVNawORse
rCDExewi6wxeeTMR+QfLvl/IXEsNymJMgzAxbus4ZR1JjMDUBNU6s3ESwR0brme7V/hmJt5cg1Jd
FgSDuBLRAVHl4Er8jB/N9aVPk6B+QZD49aWl+lmLzmt2RJMqIPPumINVChYoQWXdxJAv45f7JwZg
EZkOekO80+2xP7FzVmjjAwP2sCxDgOhadJqAJnFrn1+VGZKKmVICH+vMiH1ANI8vo29W/XZ0VdLD
5rj/qLAOpv3OYPPPulrpdiHHiRyWlWisdWx/NXLNkhF/BOcqc0/DOiLPl5FAV1hhMKdZjeoq2shJ
7XE1K+EeKphnhN3ujQZY9gf9uPZEGD0i9MLoHWjVNcXD1ys7d31/O5IGjn+7+hAV8tT6iIIyuWfY
pGm2M2El8fRzyiPa0XzvvfCwo3tIAjwSwTmlTXV4EhU9yIcLajEzqCV+o78Flf7blK467MjmZD2w
4S3Frng/7V34ClGSBJ+Ze9PW1r+UQOPhG0FolhvBby1EtDPMmhPd61d0PXjqwuevcM5s9EZ2b8MY
JyGXxro+Z8kWB9i6STTg4UGqp0fO5x+2GMoWBuyZu9fzsXsLdkO2V9rsXDWw+Vm68nY4OGxZOi3O
p0VjkwFZaWPNpczKNRQ90HYEaNPEP5NM+XSD1oo4Hu8iq6b9JKbGDVHqF3aav+W6Zzv/Ssqfeb8m
uUKyCbisyyvY2pVm7A1jFXYyNoNEaqCZIuoIt8Go0Zu3CjxOq4lQu4u7pyhLhHF2AbrUsr7IyquO
Wy6VP/cXInDxagS/UdcIJYTTOl1RQIX2q77xlIDO34j7hwBwElmHxUmJuCtZq+5bpybJWkuBUFN9
5fAvlvS7IFuoc7n4Q20tVli8czf2o/GrUkgncocRFA8bupaZ1SbKxMMRCSpUbefuIUOIuXFNXcR2
4eKxVpYcgWqmS6fbi9V11nPJZz5xRfgaeLdg7cPBiSxbls5dxImeFl8pXm9UZ09eBl0HteqH6SyR
XdX/31A+fXI12udUN8gWr/zcYCF0rRXWnxwlx4fOZZimaYlSpw2ChzU7OauKc58jTs0dp510aw9V
7R1yZEk+ZqzgfWqXxJ9m6CrA3U3KaUOBZxlOUptWd356HXwvZHVXXIGh2FeGAZyjsInGZHOKMYvZ
KITZ+Q6mOxy4fx1sHP67XD+7UgjS75AgmyfKSwtIa3rzJb2CBVnLw2NmWNPxTlFtiNoY8bbrxEjO
SD0wp1tbbgKVDrhWWcmCG5PDNdbVwQ+Fkl237DMuVBIiOhRG34LS9Zm0M0DndYlSLaIBFX8Ba6wB
C6MyE9FXawq+OtXxM+7qJEJDhb+yXQGjFMk1pE5oyXkZYuOZqPtHP8NmYmfl1468edwdcyTUeFdI
JLwGwpE8oOspDgreaUfrD++P4BPqm+FvRwsDLLJUJnC6amm+Hf0Yze2axEeeAetbKgxy+eqoU5pY
C1np1sVUqSTVc07ORu3WTgqcQgasJNGxSs/OCom6ImsJg9A1tHjiFeEg5TBUscLkuaSuO8REE5+D
npWvcy2wrRGGPkf0HXg0TZtDTjCm7Ebdqi85SYdZ5NEYRl6QNebz4Ml/2ubk03bKnUh3xr3lhwyG
l8cHqq6zj8GNtzjJu3HljRjRlI8iNXz/wS3P3mq9DTUrXgkzClWVB53xiLFU8GE1JTYxjF6sJO2u
z349xpXzwdf3RCIOUnQjwfuZk60sptla94xcWPyH737/qQ2jFvuBkMe2OacpTo7HdMfVXm8UrpfW
KMROiuX3xy5RZseu9GUQANqYvk6FrELAv3qoVrqEbWlEkGibk3Zw7SRlFZbzyaCTyamUkOD+ffZY
yUmoljYy28/niaY+NFPxegwEa7e3SvQtTqegoy/HZyTt3/w1AHQySKv29q4IBSAOAGNV3piEKJ3I
9GeFW7cy3MDEb5d0fSCx08txqhxps2u+7CjDcKtbxkfKO+j0fUbGI9NFTean5y2aQam5O+s/hdVo
mQ4s7sRg+2VBSwK8sIYLJ6JWao7WMdhxbJ+Ck9Rydrvmo36sHfhoJ1A2/Kr27uy9SQDNb3xai3uH
C/ToweBQJRvZxo1SnLqZx25aLUf65Jc82uHj/0Vi+8KnUz6r86WMLflm/FX8QxtsY+9buoUZK5eN
yIEEqioA9sZUygdGudwfTARs7QAfYqUdFmRvYySW3hjPoqBSNuh+l4cfHlzXd8opgnx+3lTjMApq
XXxlCouEMP7fPVkaWIfOy0i6j3cPs7HsFZqcHJol3M/CyR9Wwjq7CbLEW0+5JU+lo6H+bSqN43TI
knsHYLQtZ3f9QADNu3GMMJ7ybLVj1TrZ82cNZYJEJt+Nj/U419wZFAAFsa6CYNTfHNclLutK1rjE
6b/IcPqYKELYSld3TQ9w8NX5RYdvUfFMDJh2/ETocjDGs0h3GJEQlJQRCrVTzOKDQcPe2l29E8Jc
8xr6L+kcJrgJOeFXxj/l2gL/QH0WqYAkLINbNo9fx/fwC8t11e4lzRbhz8nHfaJjekNV39fzU73o
3z+AnfRKE+ZcU75FVQuOcoFjynddxtZ/pdB0BpsK+trpk+CxsBw6ES+rXCKlj5hGSpN1jXpssxod
FOlcJKlg3i8MhiqVjQZQL6aU88kRt9G2t3BV6e3y7udZPfIq6BDQw4MUm+yrcsPVssKl+024h26u
dgIxg8c0zAPLaxGzeWITgoBV7h8Xr50U7QWPdjBt2VICKwZ8Re8TKa6qukaVgtJrp3beDqe0au24
ajaTNpT4VrP0KF6T8kd8uZC071Ri7+mloe4KECCqR+UoOmkIYVcsITSHb1F9rGNMZylkFJ32uz2k
CJN4qnPw3/FlxLUs5vk9J1PE0ZEHCQA3GCH9z0/+tjuzpIKqlHW1HOT3+q1HEIy29yIl2Fucnifk
D4YJlYesxUnFLNfeOqmbLqu9w+/Bl56zDaMZgwFlkTQL/5RQ1C5c9/UhQ757MseasRYkRi2zqTad
F1AgANUDErc3gWIZWgi1WkeBCHuBAeto9anC2JFGKrTw3QS+lIh7W8aYIq8gWo4Gsrmj9KJIJccG
SKmk18pT2ojCNIvBPvdks3/ig5qdmQytjb68mJ39HsP1quxUnrwUZCC1MJZO26XhtIDkW/9zP16U
82MMxUShcKeqJubCiUa1rFbT1HZpgTuWJlrr9GIq/nEtWIoSgc2yiZwBoGKrxnoAzY5KJyKIlIKs
t/p9AEmqQLM1vdxwuIVIUExuJI2YNY0ZyLd5Tsq1eO0iRE5THVwAz11K/KiDUETyFVg3FDMAJ8kK
zt5z5G5FBD7Ci32jBthG98nNOKskMGtysTJSuW1NShjYn9bQ+eFgLyRJzE3IKtA6FDachNsPrC44
IxNWMf4HLgF6x05Jptt44Ax8pGLpyyT/GGGQdANhhE6yxilaESuJ3r9H+c9k+ZlyjDPck4a6t6mf
DbwrgISd3KNVeycfjkaqRYaXuHThY7P6Z6ri9YiE+yLAy53nATfauc85o9YoW6xuWeu20k5t8DtB
p8gZspcgvdbBnZJZyLBUjacnCfmLswVH2BDo3T7iwLSVIz94HvQfTXdWiHJfaLsnpkfYysOPAK2+
5/mnMfDMRGtm4v+3VZ9R7RrY3uFt7ZWGnoBXPrv5X/pMoD7KMNHs1iGazEEcL6HcXgRFb7Yane3r
HtgVdo2r0SYzuDodqNsfbL4KG1wM5XklOg8s5XbHprBa2uSu951hLM2kIUoI02U+USSkv/HycykW
L2jFXVH2UDwQp7uetVbli8iIej2OV5XptG7ci82pkOAC36o4+94i2LKaeZgFnQHMz0v5/tnKC/NS
/U14IAsyaHIAXNaESomge3ewSfDWvKB/dx0pY72uKhgP8Z/OokGBi4qcs/SVCdBw2hRXD9TlE/iX
ebVhwXLRddCRpxob53e7JtvJivRdjI242mwr0Vk9e4SR5Mvmm+g2kbPnl7rvI3Z8rmt6w9qTQcP4
HtAqSdFuwY4lI/lrtdsytiIIN+3CwjFhGc0dUQeO3VpXcuCyMv0oFzZUZ6hwBfyXa1oZ1tcJy9N/
2ey/dkHLAEciShRzLNzDUenEwnjeX3tI73TQMUrM3w+3WyvG6IqA6X1nl/c9rPJFNXzyq13w0/eQ
Kc9ktL8EGbGnO/DAOzy0jwollnx2LSJlib9bPZpBQinkf25ZNeeuQYyR4Nm7HXITtFF+V3+PK3c7
Ewg0gpmu30haAqB2EK+0mrfMfGbPy5Qrak0kDEh/K4lNjQbcO9p9MDeNVhU/GNffUCLi7r1ai0xX
P3VGQdNiJA+iezUCtuJhCV5bnLn2zaujhOaM5P/LgcROradMoG70K7beoG/UbtgP1y0/I8SN+LdM
rkOD1Ner3lIZMuQbdBXzcn1kAhoU4narcLu5g+xVA09iNo16BLg/8TXqNchA3AhZyTqBU0GtnKX+
ozZIK0pRrllWYJXtqC6dkmTrjZ5+b7cSJjG7rDtT0uI4OvpQGRlsnsYzX0juXq/PQ92Uha1b1rK+
YW8C2jqU90WK557DS2f7Qs1IoOmwfnIVUDZBBXI0gdnTa7gO4/ecxyglCsnt4sTtXWdmDjfEOGVb
oedgXsdUJxdZl3BT6j7OhfzwqNeLQhbFL/Fy6nYAbtYO5bQbU7TVrN7gXc887lQGuGhK5PUpXgPe
8cVO8xWZHkAA0wEa22O2v28J1onqd2R1UN6a7H5djRNeO4ZfQcg9tm6WpsOJ5JsTH0iAPkCYBoUx
lOiJ6TWtzPUay//dIZh2g33lCgwfGWR8U8miR3HOnv5oR1HoGhoKsqWWw+sLM+bgMaclxUkqZcpE
1cvRNVWHq5/rX3K7LrPCNtP0f8GCUxsUvRcx/TGMh/Wzey8PHF4e3MHNLiXbw3z6/YW/c2SyGCJX
4wCsMo6rEWn+JmhypDDdjlw/3aw1q5QCrW8WYZl7xhU7tDdd3R82jXRY03BFOvkUken2bNp0Y6aw
W8Wqu3Y+OqG2XRpnGUw5XTKJlVthOd7WztBUGAtTzebHRiT0+mMC6Usv5b3eebYjLgJ75f2HszN5
CWbn12qPvDpRtTYVUPDeLyL6v/veteopLzoqvUAA2/FbwUOrPyId78j+a9OuwFlmy6bLXWUJG0Fr
uxWtETo35d3gzf238FEa+nXIw276KbP0x69T2rqtdKhVji1bjk7ztMiRfDe7594zcfVrQ+AarOPm
M01I9IYk2WBu2s0QwfuJqy1XTovDneVj7UxRLkbIgiayOe2LzYR7UPAGCahikucMXbLaSe+q70mV
pGZwoVyFuoaMr7MudzoqfNKCbVOSnmc4xwqvvcCA0GCpW/GqPVDjbd+mn830PKkcx/GvBXlzkp8d
KF/ewMUvOFXcppAvMxbTJtLo/KcDQy3nhSigpCE4HQf4Q8b6FIc8ZUZ8XdWCuQGJGlxEezTYd7xc
SBJvMf3zDn5+bdfCC3xnEgX9OQ9cDNcW0crgBWqea+laYtN2KhvUG1NgXnnRJ8iTDsVGK9o17k2e
UrhZf6a/2L/abtPHF8GjkcSUsNrub+2DE8GO4DIKLgnZ+sXcaz5/Rf3UGRR42NUxpYielunxx1Hp
baQLnr+y8GGS65bRMFVC9gGai2/Nm4lRoYHSOsoKDuwFKqr2dMCFaWCj0lupNOaVrsXjhu86fidK
ESQ4JZlHDCZT6KnL94pqPTc4hgg3R5PMbx1pXAAolumFuWi+7nkawbddbRcXtUcK/Lqy0OwCtRpZ
IJo2ght+K8Rp3teuOLwiXG8H++lwGPWTiEqd37E9fdTf750WLvCIjvJeFDx+wEAykfKpsEifCKE8
Lq5zr28wp6kQO2jzc/wJGwT19jX5dhR5+k62tUK3ACQdT/1+pAjR32svb85oZ3fnTUdjA7v9efgs
SNxLr2mvX9AJEqD18MWFNBpfq38RWIhcmp0LacJg+UJkF86FN+0wbkgmxBD0IyY1FJIYVcHOcdaG
bwEaUNRvrE1Y7vZoiyjQexKbUNYM7FAavmqcKphvDp72xoLnjU75GXRkJhroS61FF3XYohB2jnl0
84NNOABGEMO2mubS8DaNeeq3rlvZiQh7dmcfg1AgIuux9CnF48rjW0tJrOMdr3mkMCCWmV5gDLYX
gXXu60N3QAYoaVd7IRdL5rPngVP43rnzWU4ut8EyPvqwZol8Ad/G9H+OaaWLqWSz/B5qOzlbU7MG
XHpWPG+4kAkjHSQoIrLl9xUukU3Ke30WqsNDyMKsaQ2hGhQCQFTnytT82CoCP5fuFTgS7MI1WrDE
3iIRCxuwatNteaAU6xaQNNQ9L5LwtiLlKl0mUWjxkIZk5olUU5yg6sNw/AcEOR8B9ojVKCV8CYnt
+t1TisBi6UXrRAadud/ynBMwMViUgtkyOUbG6u0xF3zr7tgJzP3NekZFTmBu5Gx4SLveKFGh0p4c
r0WDQ2ebjN+P0NochkwB0pJkL0K0v4Qq5jpUxdX8onrq4lieA5EZKObzk04botmvSuOxUcRCmv8h
SfiR01SNqs3Fr4h/rBDwXvo5ukRXcZZEzqt00J0w9DtYZfKX9ec61DOH//nJuKb2YmiUw9B8MZ56
K1cBoSQ/khJNulnIG3E7by3hRpUlhPKjz1QBjQGYRNXFvf0bXuhCNzUb+jSjQ7MlXF56SWrnxt1+
iatJ8TiyExHn4uV9sdiZSEMNrsVeVI+iDWsl6oHdFWZrE6XE84hsqAQIL/+akF1298tOsX5OWRgB
+YqVNLvtZbhY46YzoiX7yX7YbjvIgNjbr8t2nOxL6Av7SVUHb9peZWWkcIx/oUYbJVigqRpDEHrp
h1U7+pS11Dg965eW1dKY+fQFCRKVRw0aiAYlczU8jR5E3TYd3mhgWfrbBqq3DvNwgQ7ExMHT1pwG
C2ZEkiAVPvrldRUfu88S2ZRlDgS7jMElW37489xjdDXN8tCLa3wpyQ9kIc6tPxizSrTnJa4nnRZc
zukmGi4AFappkVvloGIIA0aWGMi9G1vQo5Ltmt3sW0nxJpbUIN+j5/Z4+WYF4AiNrTOTcJuYmRXO
nMoJmfwOkNtJo/B2hBrK5J+G0DSMRpigUCbf/b1L5VZgUQMFi+LqiacEVTh1vduHcNbl9qNcCrNs
bkY27zNtKGbI82ovW7pabpxLy9NTfORCDE35OV2n36Gy8RyhP/8hAkS52GduiLi2zzc3mEtl7xkI
+s0lMMkBugvCxtjiuueC8lBqqNvwLau8prvcBdDjPQ13lj7ukZQwFwnYP1vG15ChCryFMTnt5Ik1
FI0iW4Je4BX/E+ftxfFi12abyO5Hae+qwTfNimRscHwMEqSxRl0ThMBB/0w3s6riyE9BZK4hrgJF
+v9VQ5v7XEZ8XdfU6yPROPxD00JhyYnpAu3CSVBVIzA7eCxm7887pkTKXDoMrsI2XaHyRWvAEsYu
rxOrS+8JuNSWHfQKfniKyut4t8hvIxEthdZw5CQh9Y2OeuawkAR5OPotXG2M7+kVpicB8Gx56z0l
SbDcMWjvDka/NngazUkbHlNVsJ0xVQvK+TWAZKbpeoe57BPDoTScO++SQm34TS7ScT0rYvWKDfx8
JhvP+xLpLyENn2VeH383Ew+wmWK/uKLr/VMMRZGr4F6W+rBbRpwtXx5Em5ok80hGAWqAwa05y5PE
iL9d6mUGPKu9fxNrYZLDVXq5CdKqWke5UiorLtiKWMeYlvNPwXWCY6LimpoAQIcDmTfqpY52H5sK
mA9tJ+JkxvPsa3amw0ttRyge2UmDT7pwm5PdtFDLk6x6MTa2ivj7t9kUe52nzbgNhjw9pikvd3Vg
n5YwUIH3UdmoTWbZeyvxQFrbaIEgTcQq9megOKcDHDWvRh4HqOhYatojfxMEQr6S2udxrjFX5Vzm
zWXxxbufe14XmlgqStTkRDzuRj6CFefPtZ5jpDjuTNw9LcOohR1pMxMdK3vDdrUapwZMdISXLHlC
HLJMeNBHJBN9ozZAz7ik5N651QZGeqsArQkMhdefz3P5bEZhfVT1L6bF6l2lS2B112tqtF86c1fy
+w9avh/qgg2mF5w6wGA6/vOJc39guBkTpTG6TPLzn2PY6Wa6m7JS9eRG+DL4n0Y+3T8DYB/l2p/0
zOKz1aBQZ1NyEP+21Y440roukIX0IIlxDq4DYCai3EK1SgbxXV5KLKSx/Lz3sUpW6+c/gZmsbp/T
DLjo6fAi9KhxP4DOd4PE7sGqkejTS8XsFT/vL2n+gavCnMoWRXWKyIKmJWE+yYjEz4sdq3uGYzPb
rBpmRVIghPCCjQymoZDkEmHLVz0BzOxrdMjTrKAUU9AMpuyoO5eR6sLulD6T+azXIKdFDuYVG/Bs
RocoooTfQvNiRtFnNJh3thJB3YjwpyXJd4OyNzoIsRlYfSZJjrF2mMzccNrKLyC85cLUcwguBA6T
1RaLMjdbxXwezhSq0NuolW/S4nhRW8zhW7zkU26BbJ3OABf22U82CEE+dgev1Tdk9RO4EGQJSrJV
09pxTR8Kof58VeEtPOyQM98J41s8I/ZRusUUBKbcGtkZWcQH8E+I83r1sreRb6k1Rxb1jwX8aylD
bZWpEel+S+F13gYUQ4Lr7GDCWYCfE/4k0jnMjlPEwpLoRaGtl7cQM3OQQeWhyeme7daNBafpdpFe
1+nVTskDI4yGKN5toMywCFEDC5mu50sPD0CVEHfWbOmhnJJ9uHLMgvZKsu3LwHp3r+02xojSLX53
ve3QeflU3d5b3cRF8j1wdddwV1C4nA5VWQkMhnOgTf4dWPr/mlYdVdZDiNEL3bUGq31bdcDgNQYC
uFjjHQzLYDP0o6Gm6Ljux9vCR7gTNRoY6ruzO1q50PHQI3ixLf8U/ZQX3WRLh5aMHGVUcUKS3juo
U0Nk9gWQIJHb+tZq8E+QQUAQsrMCKxcAKbDFqpQf8wu6eL9sp4pkV68NHJLmgbsxJEt1aYcEA5RN
GPZoCZ985K9reT8obdrF1Zdx9V6i7aIRApgVIWIzQPDf2IF8t97Z+nntklHMpfe4drhFxI3r0YRL
V+39t5x62wsx2lmGu/1UyWakYFX68lrjP7j5rxUBPuGBUHLmFFcRKVc4WShAf5uRnBlb5NkW1iMO
F6S2l6A2qjaKGnXIyG11PSDMH7R1mN65RzW6Q7jCB00J8LR37vo2KURDF0re5j5FtKOFTwROfjnf
Dh5ea6fKKnTFhvns297AmQ+9ZKVeG7qjRIzglK6zgweIDK1kCm4WWw3HuGnGhvUP72RREM1Pg6fd
maKOk8sVx7De4B0heyK8MQNvtKCHPZUK9pd5pU7BE70kCKPFW07GEeGmBuqCKu4AZQe+nF66pmZy
D2snvqL68dLMEcmGMX12MkX+plxRlDEsYLrAWWTf8KTVFdd+gDC6n7swsJlpeSFhQhWj3iYjeKD8
cTlOjq5+EmJ2leanSO8zY75EOANcZgqSQbXqsuKaeDcxabVcQERZfZ4cXGGUJf2ESKiHTevEwG/Z
aDVRt+Niqy1VWtEeoLtYys6cDh+U88eNwvzZFsigfPymhSsjvKFxU23oJz8K43Q6WGHezL5xzWJI
hRzxOC+aN3nzueKMlIYMrzedlY4jo3oeh6b7ZUeQTF3Qq9WGyogXcM7x8nu4x50XXo+8wZox5yaM
GC6AnDRYVAURJaMX87CAHX+A/i7ON1QoTDVTbda/Jx5DRuLrfvSuIKFKltOUVZi38rpIe1PMdS+6
e7yz5hLp2IPRaQ9HselWvQb3R63cNJzQr79K5jbVwzswlxzZr0vN7buNliFc5kox2GbTs+HJHokg
O8zZpEPo8HqdF/spzc1kkcDyMXCovarecCl7a2zB8a/tyPUMXourP/rJoxm+FA2wDaGIIO30Si6e
+lr61WHrdz+S68m4XHRwnTLQ/1zV9mje3GVQRKNi8TT0tSZcHCreRj8By6h3nfi089U7TYnw6jk3
3D0gPwOWr8yMLJt13KH0wOuMNS9u5v5r0m6RjWn3lIrGpmw2OQwjEtM26/GUU/mw7VFGAjzcKtW4
H8jr5B19B0+URMMiDPbg/wFVcu9NsAHFcUrIbme6OOUaKFjJNG6k1MzF8xnUaxqUotjQ7GVhlOQL
/zgOYQxX1b5uDetLgalPe/bWBo2dYs2QLi4qKIPdWQqfJiYCEacC8LHsYA0tTDUq/Gq9o8I/OX1D
BM9dzCEDrMaGxWGrlCCkM4DmF7dyuFkVcyC0r3SrLyQOLUiDGs51nIWVLR2F824dng6QItQJ1Bh5
AJ3NSxxNWhOj5hr9kzYw0hHjjOsT+ZbakofcGRBl6BiZ7Vjjir0M0jnkd8X1LuRA+BSaKYAVy2Iv
pNkl/GOHiG0wIc9jC0mzhq43Zy86TmZxuN+xxpKZrofujG3RgJyeuov3tc1oeG0D0Ao+rtBWA2im
2A3RgYM+DNTA2HR8ma4e5OCu8zye/Q5ZtvBJkI6MZe6409uQOMDDkUj9FwLKtxon9i5Ec92OvXoQ
flECi7+Lb0PLyIgitKafqKct7IZrs3ewXWhuX0ejY2P4XwS1eJdAYmzdc9sYfuPDcGoxNjYwVSLC
agdwBGFQVo71IYPsgKa2JbdBIIfg6AwjQ6aZzorD6al5XoY6RCP0bLMKGCRAa13L9SZ4Z0qW/dJE
KNrWns2DuefRFPaP/BK5YVVx+S2uKrh4hVd0KTn/we3n2mGaz31X7n8htBYwxoMLCc5kg1VOA7fH
uD5kUcFxnq/Lszhs5lwMwuIY7PROFRGYWG2nDN4di7jSp7DSaZ+r7mDKtKJVc30j1T4MP3WeMlae
Cr6P+BQ9SoYVjEJuI0SHB/HyZLwgra0BivfMr+doy+C06WlPKU9xbjpksWcl70DxZ9/wx5u50eMt
B2BB5QldPTTZ/t6I6bKaEmytV08eyw8mSNdJVoULJyoqD3oWMFE0N3kZBvDkg2F0OmKaMihFpP9P
gJmzp40mUl11eh0ZO9Btb63aAvc0cQoI+h9DC4rMAjlY2PvaGCXXsrAxYLh3qbQWf9YAHhiKhZfT
xYFsuNPzXJ1HZubsTMRW/S0vaxTa0By09J6C6+xDEDPKqnARKf7+8eSPKhiBI+j5CoEVEoKOad49
PyDBBtj5byas9+KViU1Y1ZaFcAxTKAxAmWRi3jzZcrMV2R3lIovL4BBNB/XtxHpeyraMVYvTxgW2
GgGrJuQYtPBY7tHihhq35uvqCEr9pxbRlKaTXOlFjV+M9+seOjSGMbyxH+WMtP75okesEh0W7fgX
2hoRcCypCA0n/s3gpn2CwRHm4tZ/KB+B5bLgY/PgSyz7J3hzjQ3nRsyq39CansGD38GSjwZnqUh3
CaEo50mV0PM4uY7kxIf0gnBSFFbAMuIYvwGp7ryZxLUVPAuIXD5kvP/wVL84TNRgz1AVG6rjs+t+
/6SLCKK0/Frxa5R9xNp2422SfO2OcL45w4WfKqI9jUREH+NvwedNB1UIZqmyyHfnKt5yBoJIMUrJ
o2zpYSQ8bIbDarX4hUsJaKBtA7WGRD15IviY/4a283lem92k/yrU+miv5R9R06L4diDmUEEcg5dI
aC9k1rmslujs3SqHH8LJs7DCscbO4c8jqS3+xIiV2KJWkbHUqKbKCIHEW3QpQbp3bDM2IftXORKg
K0gHRn+EQ0P0NEmQ5F7a956+w2WNR+qoDEr4WMxge8LxY6E+xHR5nhAIivyRlXIdV44UFQij4ZNE
MFTEi5Y0uo6patkN84+xJCsMx1FzxCNqfvwC7Q0Bjg6nkHZYOWRBmN+C+A4J9JLRE+Jmn/0H1PZY
djhCFAF9FgcHJ6mjs9c6O5H9+DZCa5LFDFfMxL8tThqFQ1aderoRhjXq/3lw+c/ms+Erq9fMhHBY
sb9/Jl9VeuYqZ1Pl9syMfLUAAt5Fz7Al6M4tEbFosbmnqq1H+sSTQW+2MlFzBJ0j/zUNpyuS5XQ9
OgD54DC/eVE7OdZ+YAasArQ7yXGtRyi1to/e8YSlhwT7bGHTEauulAdpeyZR7ZTS8p1B1VIAn7EF
qfr42sHGOSPXP28wYyMZXKaEnD+O/+ZSSZtG3EZZotaAAOsPjX0tJElkr6CjC+tTH4/W0p5ML+m0
u4k206IndUzFvTm45zyUKR6wRuucZ40oyogU0ZLBSIr3qsmY20OgNsFxlaQ/X5QFzJqyC3J2fRPA
wiMfK2drGTlNF49go35NqaANrsbjzL6Zu3gpvwe3efONMRfTtaAL3YzEf+1dcOQzMo7jmFJYt1Zp
9k9G+M5eWfM9Dcwisw6EuvjAh4BUi30P34yU8hfj//hwMRwlsinSnH4woesP6BtEDjvgJYwTRFos
38P3UXCisnHatVyTm0q4ccHida2jTlRlxkY8V9M/d4NJSlW2tG8dV4fiW6ObetNevPdIpmBt3NHE
jRfVKEI2gI9ma4DB6bW5Z4yN29NrwzNLyLUBCo8393ggcEyVW/I4w02LXI6r6/knsDmO67+nEZw0
wG1odciRn+AREKI6aEzKPO2qO4O94/Xqrux0JX1zC/BxsjkESt63dcvhixSUMBTt7ueYkGLV0LHh
HY85T1URQda5XaqcSmdi1NJsZvJNYams94PdnPueEYdgHrqD9y217rAJORLKKySt8bkddOjR4V5b
MBticF/M9TA4x03a7guZUFPulG87V3VtpcgZXoMYKuGsdNSGoQ2DX/2lkHameq2uMOPzRF5ABrQR
tqTDlooDyDxRE3qcrL/IRwRsCmDTu0CJVrpbJXiRwNGQMQ5wYchFDn7zdRXontJ6GfGt87ES4cfr
6sfv4aTHCdtH+H+ctT1jeoth8kQzW4/Jn0Uia5Q14h6jbS11QRuGfZwllmpyBwM3rgJ6gww8SEUV
K5UbFmy99g/gNIjebKSZb462oRfJyga7ls1FeSsdIqn60W5ZdLCNLGsJdNaS3qy5vlILQ5yRdwyG
jzyi3U0PudwTREQ4ieziDFpG4MedU9hsabTrJ3x06ysjhTK+6R7bzYkLm99LCM+7Nm5Zml5Guxoj
xa/LWyWjfTjtfBszL1AimWIsRNo/KNDVcfDlUXbSbdoRfa+WPkZ+E7Ob4rhgk0swUDWvLd/Ph4Va
kTFfIwvSvjXxmyg8kAtYb3LPEDMltVMJqmgCJWEkUxk8zXDa4tU0wECUk87A8rnAcmQGf/udEc7U
hpzkS/qRQfK4M8fl79PjQuSAoxe/uHEBcBypTqLyD6e01RA57wYmfXwHIrbAE7KSnoNOFSQyRkki
tpE/9VdD8xDwbN5gdQI675yZtkIzRdAXIl4KLljK9oAarVkwFGO2KbY0gBxcPwJhUhea1gsjqSKy
JKOHZlFrrWMxvxSaIa7wjCMPwP8FU4rRt66o+OZQHeg9qFbB59bjVr+aaTKZlLRihCyXvnfAoW03
U2zTk1IQOMd/eNkHwWfYnUSjoLoMkWLGSSkBDb75VxpPG0wK3+22D93A1dnTR/KtEiVKEPGdUper
v3w79Rsip4gdCisnjDa6szNyuWoN8QYyT4lFxNBAQMg7BE8+NbrUjFcrvIwA9Xt0l5E6zl8b22YO
lrkBS4QJ9CQz8FdVCNJDrA1QzpBYQP30SJ6lJ02+XOg1JCOZekpJtgz3H3pbZALGOHSCwSziozPb
cR7eSF/xwDBSDET7Q9T3lmmFOJ/NSKTkTv+XM6v6FTwlllfyjYdljA+myg23DMVdQdDwdqDz0Xgm
7VKcJrgn/i93q7w26GvT7JVLaJGK9CWIUoLnGlyRIH833MGnU88rtmjkMDEVeBFLJoL8ezY0rfZT
K/ORxuqcyh8I7hSxvUAHHwtE82+4OnUuiyv6M76G68dRHboH8eE/BGEkLYe5czNyP8tvAv46UHpA
l5nXknvoMp57c3s/b2AMT/ifQthrLhnO6CSqSYKwkWg012zrWYItRREWRRxAMTCG5WEYHAfJoRv2
eOIEtIuJHbvbwhiPUO1sNQtchOw7zQihaAn14hxnk1P9VDeTS5Ghz1PpZH1uYSGu2+q4NFhXl92y
Md/7ws0nOAtloKHdtTSTmn6vQ8EpZqiE/6YkoNhtyeQi34z37llgjFQk6UVWLmS3Y9Un1vq0tlWj
M2SxtUJOGBON9By5Za/uaRtUjYpelGVbHGyUbcP7WwauOYT8X9l8eCuCRdgh95mFfTFhXs6bu+ny
Wn7UbiakntKlFb2FIocV980dopWHRmaBUlSr5/wHIt2XdJV13PJ2r3Ff2atJukm4bA1ITRxXw1ek
R008INvZvYFiTpCC2bxqnQPCVwmJkEIszwySHElJJcVvoBVyNb+Kf1c2Jb3uesRbwgPYV1yHEXOo
vhTjyzvFJdaxLh4YWvpmTxcCn7+rV5LYCIo7JtMWDeDM/qa3XtfQiQjOGUY4/0iuOBoZNppKyUk/
9v01Pms1Nmz78ZOs/ORVAfTLb/hIfbDwT619cgoG7gqn6IWY4x4kljvrB2ccRBWDc3rntKD637v/
jlnK4vc5nKKDsQ0EHLjrAxZAv6r/X+UIRRBIJHnlWK8n7HVFpP+W4ZKaqEf91OtjTm1C0ubQa3za
+/DNx+noGUo/Q25Q2KvTSEB0/kxZD7E6ZSjNZ2o79UEEZ1Zfv4n0HkprcDqcA24CjazfbZEQD5t1
yMpLogbpmqi4djotzqwmqPjSHyWxZR1ZpPXJ1v+LrzpYzk4fg0U9oowb5zr7bpeLdBaNECaraTHO
SEVnqMtPWEUV4Cs7Lq54/8VwLyjekR7NMNyNJ+fUWxZNECe8ap0PMj0xZfhoFjgHP4ff8LOYEHqh
yOv9JgInVOlDuXlClTcRMIXzgKPTpjQLyWhFYuc7JWqtIzvtoIIjq0HeNe6KuDx0KwfIllUkiKqD
Q8fHo0ZqHn6XBAy+eNS1/Nlsp7/kvEpQwanRY3C9R0a/glgDHVf9f8sCoGi8gRm5w/VKgp2RnT83
L+KaOszkr5J1Z9hRVls2vLC3Db1Nmmm//qIphd1MJu0RiOP3vawpjlsDYZ9KhhObGIUtY6TvyWzh
UJnc5scs0o6cJvJpw+EXzEONH+M9TSsJyZjfNfe74XxgMYK2F//pybN4ISPH9eKFOujDo/XkMSxU
XrQYFZZkvY98Kda8iVq4VMPJHjUk/7tdpRL18bPERYLTgSpcep4u42socz+A843ueXYdsvTzKjyv
GFnQlRD1nCKFLIrWNaNJCobzF28MQQ/ztVVQuWEMpY+eFKwj4uxQQIaQeQ5FliVYurH2W216R5oV
n47BP2W7Vr5OBMzfmcuRL0u3AoXqWRpqLT+LtaYg/z4sT8D7GL1xx+eiGKOwi7QcJHlsfaq97yLF
yEZh+0x8uRo1EkVGiutbqPuplXw3Rgvxd3FLhb5B7WZU6rVcblS4vr7mm3IarxMWcm1Y4qBi7PcJ
eLfhW7NZkukACig621fJkqNirYbp4qIZ1jnnF6tcFoemBTRUpAXCBDqewECttZPZjYnJSECEbqTc
xgH5/egf0mmKwoeZfrdMVxrgGTEHWIPceDYGoJaQCXA59Tc55ZjQxEohwK7CuP36MLSspPuA2jtO
VH23nW4dARb23Fd4nh4dJiuoe933z6Lwpe0enAheiIiZxvKbDvVNmh2W48WdGG5y19jyTpVPW8hT
ArS/Ec0Kt29lwyZylC6XVM51BsZneOXvZOdOjbwPIekDsJLuIA/WIpXt8DH+86LoOCXBqr788Aqt
Mvo45fCV/497yc7ErwQ/D4BdO7s9oJ3l1pr7E164g2faziHokTJ1a3rMK9MLj72gBhN1SJ48PexY
WvN9G9WwnnZkRFuhXDO2vzNJnOlYSevx+41SfiE5FhxGqfU+0+Adk9VMvVUW5CykdG36nknKvG8G
+GPCubvAhkan8lyGWIZ21N1ujDk0Qtc/1U6t7OBbkSPQd7azvwEg1jT+HA8DNeFqF7LmFUYP+q2X
00CvIlDhxWU+shD5vzccTcHroIWTCPLOZdrrhqXBSky5fPRX3uoBD5qkTvYo3pOYX3NfvdrVVP1a
ICkWOsl3NZc68++Vh79LXkuNx6TpMW537g0zNWBiETa1Koc4w9WcIi2cswRiejMCACw+asQ4uQRJ
ZFk9BWlzwkfoH2psFUg/9fxogkRQMc3i7w8byiDQZY0G31m6QFdrOkzdWvwOLGQUpIWP1BJda53r
nz0dhWsAwireZl4td+6aS0xDkBvcmZyN+6mA1BCxs1a68YFZbhlc+mtOrO89CFi6p+GAp5B0tymC
/lDbmkCh40ZqA0leDQyOIvPh4c9tr2yQZau9Ois3015DAuX+Gc4LyycAFD9m9LpDAySdjRdpfTsR
O3J/IgUxgYxnsj5LidoqhEUF1xwv3AJ9391Qz0cm339M2QsP7HtqFYBKy5HC9/OYOhwjleEl+fGx
0pWK97Hy6wS4sakGcpZCOl0xY8hx0cZyvNZVD474bQGUyn9BbcTXe4ZaiO0uN8h+gRtTCF9a/62D
SApbHcVE7xJuMBA5KqUoej7xzI3KmydCkGazYb4TZ7zL3tcUVo+KylKDZTbX53KvKun0GwVjmGBX
jzFUrSvTufS8vyeWiEVriiWvCAGy0qp2SJgtJlhflZj1pEjHJGKVsSiFibjhRMuZ6JXHFrtbMABo
lzC9k+UUwkkZXV+/e6hy7BpATOXr8/aKBe28I5eaJfsr32Kagz4qmeNI340sUMykJTMjpB6A6/qZ
R02t6dYm7IQwJIEZ8bg4+4DXdOZX7Mo1YD5jGjwK4wXDwae/fcSCLi0y3BwhZzD+E4txBhyLx1Fg
gFqNnrgsAWZPTgJhz3wYIHynSLOBSnTUOwUhFiipO6rP2xJECLPITlU93TGW2l+x2742sf3VD15v
CYvkT6dn1ZjCCNDxEzXpR4On2u0jwWypukypa3ABXby8U7/D1GKgM2KYrZ9IR3IpWqd28OINgUpY
TQ4PHPcPUUsllVGfW/lQigfx+iX2OZ5ichYOwo5c18V5pkhIGKnVXRBChPzJuPFH8RcRFeBx3B5K
NZrmhKXjGDMczC/Dq1gq16+aP1AS7h+1qnjYO0gMrhY+Ny22EYeJdOmhHU+rvb9ii4xuB2WGFGlU
+7FJvJ29iHz3OG2GCHMfcc9+/CNimC3IV4U5rqhnKRf+NJwBXIxKvLlyis6tT0mNQ3urwfyeQzBB
CHoUtze0b+DD+mxB7qntWwg4jk1iwiAg8sqvsYGIz3qA4v06vB+l60UTWhYsYN7m3QBiL8GXDoWQ
o6kvJYkD7S1mzNTpi8D95C6cLU9I6l0H0qDneRkF6xcB1PD87fYzZ/VJGL84SmT9AYWLUEThJ2kj
PfXUy83Jfbjt/iabPnO2OvWS5aEshQFTbFkBwYpup9xSI+kVCNtf7praB/0IfBP0RcPUIJ8yWaVr
XRuxJrbUZb4UQvbCkqcrVEHijLlLmvsIYcOFEJlgmEMOUyHlo1iWIB2eV2OZJtBlJKH9XF1d+49m
ORtqGZGNo3UhJMGOcM+nDPhHYC5QS3/MVNkVapEhyO2MDU3ekVlmb48QOedjxcKBxbCw0M1V33Sf
BVoWyPgHPFkV9qizDy1F0/rGl/7i5qMev5k3Ry1kstDgnmFjlGp0zZgtONXF0T+xZRqhoVM+UbU4
DEEU4nYWlyTy7kMeA0EC/sB9ODP/iY4PMO5lcghATh2v/+5546F+FdHyqzwpRJKlxJuR+2RVAuHl
VospI0y7koHzxCDQsyUj8GGQeJllvZrYDHtJSmyTyXNwtUo2O75cdlJonNiMq8rCDCR2HZ+W9B23
UCDNb9+gybX2AGAr2smZudznCIRblDyUcXrkG0TWxPKX3VVm6bxqPZJ6HRMJNQa2uV6/PujwJ5Ww
UaT1DNMQC092rT54LRlqkKpd81tSW2Y7hbUhS8ruK1Ij48m7usEwz4YsFkSUgG0PJHmheUlNBy74
jOKteQbpEF7kzCQozCm4jfNPpVfnrmCGOCGDxg5Kpgr5TEwJBlQjbOaxZdib/m9q7VdtrRIVCFu6
a8/l+Bq3kHvZywAYZ3rcwSozapaw0wl+fXxNB2nCIMAeqoo/xAKsbcmOrQoYtD0Lxw82x5bEOap0
ADw571pKLSRGWwugs5Dg8Iqvb48MOBBt3IcPQx+jWP1gJkFuejy4UvwRyi3/07/degOBwinkfilK
F76cwDGeYL+QJo6o1gl7oLrzZrxjv9E+ChRnZfOEaijMX+ESTikIPcV80JUazFPud9/C6P9ANh1J
veqxllvqBv8dYoMx3iVX3adhcx1l+DxODB6ZOdZyH50bszQ5ijmfigrdAgEq+AsWeymmeo3r9zC1
VSZAxA8BeF5Q2PCk0y0/S6QRSXQl409oYkQ/C7XVYiGqv6g4Eif0Q0NJ2PN5BiRX9Ubr3XlIBfnt
lKPzq8YeTIJ3L5WG2zvPHVHAU+kMCYLbpBDMPE9wz3Kgo6akuv7BNwaH/mnXziPi+Ra4uWWYVMAL
OA7zdB4qvRktQH9NaQV/EUWFcp8Ga+762yvMXCAAHhFlWN423Qf9QuvE5hRIksBCsNAlmHeL5Vma
/roRhyYAXuykCqXdjuV/VP7SWCsu/NOmzKJOIwa9FA0D8iz7M9ttXcXkTab5bIQJkjUAFvgNwoLb
wHnGbTaJzZs8fPtj7UkaqmtDYJbXZc8RGQ+ceqpdEHAFjNTHhD3VEv04Gw5yEYmWC3+Fadne4FC/
MEsKBfRiWjm30CYopaGzYbWrOeLmB0mFajiNc/k2ndu7dxf65x4N1j3E0SOwkiG7dBZIl/uFtu2P
E+T/MBp3tvGxYmkDp7m9vZkxizXvMzI6CwWEL5ZGHvQE/wqINJHkYEUr+NIBJPvk6HKcn6RNAKbW
aPfBfvTxi/NZ8yhfKWzSRetPaf9QCDGI18CQgFTXdLOBEeQoOCo2fReMH1FCWORZA3VBCv1eTnjK
6w7XO5u0qH2xcN54TCfa6tF++fZQAaR6ZinSrHQpMBgNQh+MDEOG6Y/iWhKhUYZaI1N6Tia34Eb1
p3xAIIzNeIdbBWVi/8pwSimaJuJTYUJdqRhtBbCx/Sr67tMUkMdl/Rwd802qtXrSw/FhZdnTLAt+
KsYwIh6apuNajXWgeVN3qTxaNEdf+XfISwjIV0NG5RQELTc3hIGBQn+Gx9UFFr8JDU35FQfs0qOC
AX5cKqxZqjRK5mI9sjOB6HvbOZeQA1o7LlgCRo808QnoBWREwfF7Ba316ezpM6JjYeZYy4cK46Bi
9vgQZtzGWSUck2UCzfO09Dr1VckgPhWShn05BWTwae7P0IsRBMYp8cD1ccyigBP9KJDLNp22cfcH
07oMB2XxNTvlny0BI775uC7FD4O8GVK+PZoGVWfaCJuzmPUVva4bCkKpEH7AMCrREPDvRXdj7agH
Byz/jatXMrHMq90c5nfAx00WQGMR++8jNJZTqr5bzMPUyDNbFVFQNDhUhlcWFy0NpaWnYiZVglmF
1VYyj2QlELzeB8QYpvZ3eJjGDR/7d8ZLDTaST0iOGF5GwEJ7ryNuJMmOjh7C9VyrkvHdCWnWfmsG
EUWpi8lOfbRh5LIq87qFvXd0HEbiYtVcQ+RhiKfRTSEyirFQU6uG2wG2YYhxfwDcbFOMzuf7sFe0
UoJsCRP1KYX4PI5JybXpdm4g9bv66/Xd0zFvxQr7j3RP4TWEhKYN/icztG8pw3NWPJc3jQEm3iq1
6xdwX5dExIoT/7QtsNzIurLQBKobPpT1a4Xm9/LmqKl3iO87W/5kHtXN4YeOtuMdUNYPdvsLOC4R
BR0uYK8PDlvv3bDHSr13wMwoolPGFN0ut9A5RYgxSsBIC2l/pvO/6WykmmOTLxquQxooRCGO7NWy
xr5n4SrA6mrqrqu4xKwrutUjKoGP3oWPVOliAXi5TrGMa3mzxpi3oDVjjzE5OK0+9p+lq2dajKsn
0kUbRWvBnooHVnVdUEmhosq1vtOc7+1/87sySuo8BvuTU/IDn1IJMW/13UK68/McmoAjBKD6G+Rf
GvXIdZTD1i7ZqVa+PiUx5ReU9tmxgmi83B3wF9lxqnHYoheTeGgKqtT6UnWEHtqtN/N8Y223VcSk
VzgWznslqYZjjjoq30o2UCjXlOuesc/gMlZSWAC+unmrxayyp8hSoiibcPfCZf93PVtznkCIWLWV
Qbyk0zRIlle3lVM68Xp8v0CCYs9AbMBNyDRzyB9+UpBER/xlOx2JkmWP1mekLFVP90UMHakFPPw/
tudsdAvdoh7lpdy7NGlpzGVHg8/gSe92xq1erMFbuepl0u96xEvCICfgluxccOh60RaNqxejRQsB
N5yekD+ARYkYJCDFP5H2vSvC1cHQm2cIrsuPZtthv0lI+lQd2GtMmbW+58Ib9aU++HErPjxb66TL
9A68qn+QmWSP7Hyeqb5R2NNxlJCk/h/re+Z3Rzc8yCljNix3j3oDKAUtQ2Q3KsAkbsyRbwysW8pV
zSJRgozukri7lShgi6v9DqPdrnLhYiqvyhsxwpA5qTmZKsoDcfgRpxcur+g4mXI7rdvNBRb8+b+B
Ac5AOgzXS3JsRYzyIDVEVL9GUEO/lXqfq/pBjNGkwrf76wMmtE+1ZaufWOUO+VTUyIa/L1dORm0N
vcfdJUk/XyOnEBA/9t1fwK6X6/C3YAeVZ+pjXuOsTQ1nlyVWoZR3MJQmhciCXCoQ33Zg/uztcc9U
smPAXmYgHraeu6LI4pUhMOj7Gqw4HEAU0KT1DP0ANw/V4oG6V+G8edyJ0Be2RBgvlaVssBYjXCf5
OgB/kotabXVylNHriv0Ct/m64FPBpWBEAY3P/4YOP6Qz92JORmKn+VBmF7b07MxYbNmq7y4bb9oa
n2GIbCovu1OCs2RN+tGdRuh+Nv1JFos7VGtahZ47Uo37CkOKnpBFvzfVf09ksQ9Dv2lYCj+XbPg1
TeP40KjSGdCMEC4LHLLbwbaEPk5qaXAZwKTotpXMF3uqgjxPyPpqrBocL2O2WexhI17tNoU73uDW
g6Fi2m8sYGCrfjbLFw6JdnTcehnd/LmFxSGpRDe/0nX/v4tVLC1Ih5KiJ5YWFApGjZfXFEQrQ43t
4wW341B1QjEo0H+3nbUkfuE1+e6A8DO8DbrBuu9axHsPHEywJNaiuNe8xk8BY7gZgN6l/D7AquB+
7X10BMqakfo8f6zQTXrK9YCvWzp93mdCTXb0b+8cLcS0DI8qbO7SzbmlrPoBrYN+i4RCrmJGVBm/
kfhL3dHAEMUm76AJSUsXHz6fWG/UwfbzIeJlMzm7hqcuZqlI32xid7zzX+IWLLCra1UsadTGzfTZ
mArtTCS2R7PZrefNjjWV001yBOpNtOBtwznsBjL6sOc3qy0zOA8puTx+vEuQ/O9ZmYJhgzYs2cpt
Bcb3g8lP8dSUGBvwuvpK0SjdBInHELRm48HXl4IdjNy3uHvzeovop+bPiMMl6Ipvuebwe3d77ppE
6i7rY69+gOEffUE9eEv6mJOejFKNornhes6uyz8kuSP20bww0vbyjAD+33Wrh159vQJ3A1SyGDB6
Aip5F/ncvhkq1PwSvobGs2qzwxur93DxsyPmQtBI8VdrD7t/2o2InVDHKkjZgTQ6VPPSPeoYjHha
jtkLR++9ozE2lWEMXDYwD97PZa2njksgGESq/7Io15+edVO+Pl5BzaWAJMnIZXGlIJFDOgbfs8c0
oZ5hq3KBXQprhS1/CWa/2mwgoPAhAurtuMqTTlbevsqSV9IeT02JGVA1Xzsn48iF6F/+xQ4hLWcZ
rfVKvtywgiqlUWT+PZ1j7NCyGHWZwU/dJrgAj9jDxewBMh7qJmszZ7ma9zStFBvcbJDecg0kGWbE
zTTlO2cVHVDQN/Ky34l/KDmBNBBxI7CU62o5Oe2iBllgKaltA9yDdKAvgmC6qZUBfwTdi0erX7ie
YXtq+qDSJN1qZrtMeGePHe5Zt7tk87nx7ZidbHMQTymdtok6KzTLeovewE0VQO8eeuhjofPRzQbz
SoRt0QbBqOabQHDNpWqxTehTwcBPFF4Lyz1qCoFrD+Hd8WTq94n4qa5rn6RTsmhD9knoLRFEGQgZ
3lnTXScSNqUk5TtvisPPPvtkuPFL6ym0s6dwHduVBCi1JioAMez5MNIk8zoPy2ubePnBFR3wMjOy
3zUeLmu/TtK8ALzPu9LEuyzNU5BzC4A3GNyOG7olVq0+jKzVCD0m+JlxR+OqiHXkkoNGCvi1YOIY
JuaH+IG5FiUHntxM+1IoruwP7CF/0YnqCXVj1QzXXm8cKXtkhyaqvuvLNuhEKJCj/2d+4j9hBy+9
MArR3SKHy2yRCCbZxJUMBrlVPzfvYn4FPJEt6enTcW+hilO1abpcvPVcEwCkB2aNevp0jFzsrwEM
BhJu2cPGmJFWiix9ixcdodU5aCMVVnZeIHCCh3utQXqKvmfYPoTT8fPoRhxJBAISuOS5peagIqva
x8gLGpP95MM0hH6bA06paltdHMZFXFOi8XOoIY5giGGXi6yNzDVrmb+i7Ii3Dvj7xatuLGdGIegD
Oopq4Q618V9VnWehfqIfdMdflrdc0iItTf7OdVrfY67bRvU3uYgpqRmUd0BiBShIbVhDspOiHj3F
7He7tVGG2cpM8f6Z7GL6Vx89uY3YmxyUK+U4W8LXd9ZKH6Ckcn6uQCqngd6knu0SXOoeNLjBmIU/
K8LLBCKlNePW9bQEim55klxeSEDoTu74BbvPWPr973yxvo0Xd5IUguUDUb/G4X103sul9bfnRSqC
NmTGwawI2hdk/VUb83VNnKDA5dakkV2Dey4tuzfI6VfJ7C3vsn0ScPoU5M93BjqWRXXQh9AezN6w
KRMeImW94TMNtJoxaX7M/1G8rfxz/b5f6tSgSy6fr5nk3xOV2Bo+EAd5lc7BHuiZ2Ix/cRgpvsOm
dhkp2ty7tss3y9OflhfD4XjUclZHcWoUnD9X+yRq5p82Io20gtAgCl8elevDEvmZLT83Yd5vcKkZ
o7aQdyOvuiFV8EIJif+r0qa1bL7AFce3zvLxjFDgECKCCed0jGmlwoL2rlcjD2nhjAdsCpK0fhMz
rk6UxT4jamM8Msf9NQnphdiW8m9gL08IuekqCEKevw1QC7W5i8qqKfmbRcvZV10+mNy+Utx+V6ZH
WL3TYhdi4FjgmeXnMzrRvCrPTvhC0NTiNdwShQkd0QdODdIGoRiEEdJkEpWV+pHdhrPTEFG3FTTm
SO3QGii2wgAb/Nv4w4oEn2xDPf/Jgo/cw05RbwqVJ4Mf4Eit+79OBoJq7rjMEWHlAFtQsJ8yFCIC
f9jGUU3sgiiPye/n9yL+qjWSt1i0HzeFiOSo2FDq+IgEuGSZEuk6vsOPAQCxsjuzpL8NvGZXIHQf
3KNe607Qa10f8WBIlhoFlrvhHLZg8esdmnCTAskWqHqdX1I513CaCJEsJHFYNflOyYTFh2bV/cE/
vucyRzh2vCWkRpaufIiAkeap24T9cm4U25xYpvu6qOUldOuvpawF0xDRajCjGDNxgdcdZHdyuSGV
jlDJwLXRiXc9PAc/dMoJgtOlElJPkudouXdts0BllKpEx0MOdDXAZzS8pUqx4TKQ1w8je1Jp6Eff
ik9wi4qjatWZcOy2uNJ3JBJExTCVmXi3OY7hA8FwhH0D7N6Z/eX49u0QHYQZGNOg2CobYdTamVz7
LaBA4+7io4i85Np7/vwAkvmdvd5hYXY+ymGFV8Ikw7fNUKidJdAuN6ki2pBlLuDl+GgCPRr2O7w0
GxXffkseInFvOtFpNWwNIC778C6GHB/WmCOIYyKwb5DcmXThI+KCfgSBlbHdrjtA2TAMDKPT9Xef
jtwVUCaQzXuI1y9VBLCt/p8tkO0vOwBPQN0S40Q0ZbllKbq4yHxZGuL4VARjpZmEXOt5P78NdcVC
djDDSdhd74BwKrTkTmwQCUxGD4igefNx+5OQg+LtOONL7UmRs07vqbxR1hYOJo7DlgbOeFoCjx9X
dEGY50i2W/ULSqDr21vaEaebvgU03+zBRAL/4eHW1fXBy6HkPPfmJBIm3nHvbk/0k2trli2N3L0j
5S81I2r6MX3YudsgQNTZyKjJgdNDhx3ONfIgxm/VdOHVM0M9QijZWqe07jNLOnetVFjrXtzT2QAp
cIvcAs2Ydr/mLXOgIQxZcUajRXl+20snaKi+3KAGaDFDhuOPyLa5EhZEjxhQJkYT5sa8cPb550Cc
nIntZ+9DpAWc47AlLoq9CNNvwcNhRxs6K5RaBDYEMvAEbgjPUbpjJJp1Jpok8ncDVY3DnL/ckYa0
xVTn+QGg4kNpRQZawuJoLeHrCfLbpx2ws2ZeZsH82xu5oV0uuQYh7FwWCr2pJt3AXJCKLh/WqSae
cot1UENSY4dNy7xo8hOCK6hOhzpb3lnHFSJClumEnSDjyWmkZZjMTQrGJpIQ5qOChujfCZyHso/t
D0HHS8Tj7dIOLnR/aWDDVgr7mvHF6XbdIR2mALTClSD8Qm/TAlSuvW00IQ6vu8rZTwty/btPPNJY
RSzLvpgxjssAnIW2/4BqQNvqaOpqdjryUuRQrLPsvuWKoFSBtP7ziiOGnH430g8PZEyRVq76Ymog
ld42GNQ2dueEkATWqCcyW9Q3+6fcWnH5mAXFdG46HvVEXQGZ8P40XF1CaKnD1/zZsSmfwND2dFAK
yivMHsdZ2U+RPcos7S8sD+TR2jIqEDp7LPA6sE+xDP61h66JsuYwl9/kq6ZFmdmiWq58lHPO7uu2
VhORfne1rjmWjQRmWB843UUZevLKGcxyOzchZlxKj4tyMwcb/60PZfYz30rR1Cc8JjfC0E712yNQ
7z7N8IuYX4yKTJX6g2OZzNpOqxNlir0zyudmLNFmw3/htYIrtLnBD/RkP7iDAVW3BOlexEf+OoVn
Knhgles03L39jkKAOimYXMPFqBI/wSr5cklvbamas6Xay6qre4ieB9lTHtolr6o8Pwh+5Fvj4NCt
Q1AcefQahJDjoWTxckWDOll3jNeybDtA+wxjISdBxCw0iqlwU3HMIfysbVmadsiyLd6qB4hezI6/
DYwEkVTxA2FJvGOZpxGLJ14vTAi9tYgrPtNSCG5MkA7s4oF47hR09kLl4Jav98o+Ryrzi/JAqarN
a6W7cOZEq68VLA4e0201p3uWaDiIp4lfLti/naBeVh1ZSdrLqOubnHTihxNb4aMznKTE1rRtGUKd
liFPGjqtm4P++mB/Aa+u7032hjhWWrGuTd9tOmxU2yFsUlv2X2+7c7WddOhgip1A0ByAJIMJJqM8
wmjj3Rew8XNgS6D1iuSVd5PaX9SuYjJvzQ1idziOx6wJharnpUZft5CwCc24U/BqSd8ppHt13DlQ
qRZDjwwCd/+ya9MfMgt13l4QHWJu1fzq7icTf73ba54F+BiR30bMG3yy7DDBSLm+KZgeII/94iq1
5s9kdntxBmKET7vvg1lBf/B+4e3hLo8gHKZAZZTis6hCfoivA56ydPLMXk/agNjSRYGJvRurvtbb
2zVzxtfUNX88C+6Ibgl0k8GSmNCxmn2VoVEjhpfYquJWEkfuGhqwYnETGd47CqGmtb8DRVn1kwbb
4RYQo44kjxDzXDRLBEplaAp9/I5GeSd9bhlkBEYfUnH5XVabKO7HkkmGg2IrwI1eFcLIR8oNuIvY
cOMfino9oev98mmTZnWfH9APqhLkuX0JxhW1xkFOGW3EKKI0sWxbT8JTr4GuYrx83wFi45+Z2KuB
wNy8/HaNbioOm8SUv6cT8s0XnWHNufImg0P9PLNDQ0ZvYVdhSi4OOSatpDUUAskS6MGjs6fgMmK5
JhvloJNBbdqMM/ifZ5rsECNCmBxaoKF07YjlqZCXfNXdiP6L+nWSJC/4gEH9bStqotL1d1EcKx9i
m/Xgc2WA3IVpAnxkd2ibm2clI4KocYucAsAE5f9vDrM2EcIJ/CR7qadF9qtw2FMj2R34vtWvwGvo
qTBIkMsXP6j4KkigH67YVZ5ldi3yQWg8YSSlmqsuykGjyudfl09yoSERXWLV4dD2NQlZnX/h8YVN
7KWBLUu47lv9fl0CZBsqF7TwoJOn2AOPVD+jiYYr/HR7vdmO+aI3QZhw4epjGIypolFOkLJaSPiZ
wfUGBn20C1vxZ7Y+MnE/U2xNdZK1bGOCvKYdReOv1icpNDDsfpV2/s94t5KHx9bH8xIj1BBHPwfL
3tLBrkU3sg1+6a/VkMnYhDXNZRHIWdpBooa/89d/AUSGZ+/r0gsS31241v2f3v1Kzd3h8yxpjm6c
5a/5NZ+fqIIZ0mj+mk0/8EPEutCFX3LW+Oh83Gy5xwMlYWe2z/swsAoZUajZX76H1uCJYWhEeP1t
rpMvjKeWsXn6JD03I7i50Mr/khJJydu2cZlGC561/BEZ1KicK2GwWI2d+gXSloTdPoeyHEvOXfIa
KDFyWTHTYOITv+goM7lrOg+iTlglQ55LKDNYUc4MCUpym0A03H9pNSgoSOhTofsvWGLCtuoiRjCy
P5eTpEdi5vLNgvEROMqI2KpZ5fQY9ms7QobtpfIZObooX1X8pG1xg0a0+ybh4N+gtnHAAabb4p1+
ZuCcW88WzgRhcMAQclORgIIkAWQI4zJa+MS7UW4bcPSFeMyWsEseoo0b8wJEoouhxiCTCUUVHM71
gS+5/OEneaV5KwDIpTNNk4byZfWexSA55HL24ThZJMUI85No/AvKPNcWqB8oVAZoX/S3kIJXmL5x
aRQbCllQwWwLlV7Nqf/sHldDH3OP81wfTTiDxASVKUcdr2HUOVh3cx125C6wjmOEQQ8esfh9WHhn
4ZK5HdoWRB4h2S4BDASXRd3l/vu+hIb2IYts07/pA2Vw0yfoLIo9X+xCFFeYvGiJvcbCezAzaxeY
BUj4nxMub9yHkOKl+yXfGS/XKg5qxAGq5bi5A5/+kWORkWiYWAzFK4v2mukwZvbqQxLebza+pE4R
IbXkto8rgRei1NUwGCyeFDIQJdH98sJ8yXUTnY3Y8UnHFzx7dZ/qq21F60CLs3WUE2t9hNWb0A2q
avlRjfLqdsiTZ7g5LW1/1B/oHsBmFFabQS3+zzWEpynYdF7qBkiThsnCVPdNl3i2NDI3lP8ZFGjf
VMAQFzRbsZ2BFkfN5rODxiXjGbggtCBtgprZSWC+yBDG/H0sOEDMFcVbOagYhpeDlWrwIPLnbR0B
2i2xXuC/XDxSWwKjGV59eWVZp8GxAr4UvDvw01q7gezzNTwI2ZEfA1DE6PUB8bMjZuTHpT14ufDp
ZZS6KtsE4F8as6/5bFjDPFWCN9uOMXrLI6N4mtqSvhBuc78fGSJFJ8bKYmrBqrcfk7QOtxTuiS4X
t09xxUFhq3XlDRQR3U1fAH2jdDReUaVdkkrhsCQfKp0e3WbHwubrsIrQGozHRpfCdkvID4uY3ZZL
d/jB3Oe/q7WL2eUBhfnadfqno+t3mF/vVaW4QVyMy3dKjnCbBCeMFr9SlvWkoJuRUe8/nIwAm6EA
XKiLve4oy/JbcXIpBS5A6KYmTDkZ+rl260db7EZU7x4tB0c+Cx5RPkft4MekK71KPFn427IfjP/3
uhYcZSi1c+MlDaTD+nT6Hn+JPPKZ1ZRxwIJmxDWavV4204M3T+MrcWuLdVfe+rdU5n1pHMimsXJw
E6xDqNLTP1jKCr0aChvVs9Qf7xAYvKtFl/ZjF7gtGDVi/DKIIcDfL41paSPxLUFp7moYAlGrnhmD
Fd2QFvd2TJpRL7GBsRijJDtRn2CQR+G5iwo0ce0tpKVpZXL986Z0IcljQXUxO4ydEnNA+DJnu4a5
cmf51GdGyjLrQKriiKAogHjMJzAHIVAuCWKTv43OHpoyl/vZKv2KAhitrMzWzu+ewHYkG/PBtt0l
GpAbiZUM796qbJLDFSPJv/n7a1O2xd9MkXJyc9mOUIL9TTwwbDgA0+cgwtTyY6TgyFGPfX+oc+Ni
kaxcB3q5ws+E3Hz4W1I1g/XTDLX8Ls58iufbq69ubb2T/MW4ICW1FAsVfSsywT7ob8auqt0hJk03
sDSdfAeHtAfhxNsHZUV2nGW7hFiVmB//QIf2WNBq0Iwc23DYt2cwcNpa7yWFQt/2tCBk3OTxDNK2
L0nCzGIcqAZmZeyKWsVs849ujZg7CRYoqLygKzktrQJOL+a6C2nldfJSZSSB54lM4aFwBrQYhfyh
R/GLV91vg81qqDWtEBCW+fK3fJy1yG/oYDERUVun072WxXWzDrGvxehsafL4NY190sbivosSRc1r
JeaiJaBMdLxTM3Y5s1G65craaf5E19kJW91UjnzOzCP0sAN49pX/+h2q35SKz7U90fTbtyl5r9D3
7Sav9g9N/f5Sgpw4JAFFaRTWc3ht5nvhbLNRzZX9+ZvIjLXDeTMXeSH/A+aiMbBmDNoKwbGF8FF/
xGh9VkpA6MqXrEzEitwRDmIjhvvIavahNuP26T9UbqT5t+TvTmetdXgk3HjCswlvN1pEfNmUHUJ7
KQhRLkkol9KxWtZkFdyzLmqqQcMqzksMdLD5rrDPusn33B2t7S161sJVzdIRB2+P4zaDTV6yww5a
pTG3ZLw0BAWH1ONl0AdwXKWmQ+6DyII660Z/hE+aT3nMWNznV7iz+GgkICVo5wWrfuTa+bHln2+v
nsVXi1XmHdoHhHFJySqlUcriYRWNDUrnAirfZeth/ZAgf50eA//WEwErE4RVcbNvZxMl0u3zoJvU
H26PYOgoVHUvtrY/IXqxlo+SxuCrIu1bAufw1F+O/gyOR1Qi3ehdBoNg1RjE2PUAgqRHh4ehWv+6
SqQA6Z/pCDxugkyAB8TNK+J5xK9SzDk/+BF8LGndYYSrRAk9a0GP/K3o0Zpx1WTsXC1e8eYpbGiq
zGQF0JZrvImT+xfmz0fFvSeRvGokv5i52gYYgQINR8lW4HIMsaG0v2TOJJEQBgEkpjOZ52NgzLeX
iBmks/QlfxJrpnugIkOUDLq9/ATuWI4ptmR2sbNwi9m6YcNmXbCzv9dM+2tlYmZ+Ohu6GPm5/fqE
HTaOyWuI5GLbYKnRPqn/O0d0vh7PPdgIrw0ppvKq6a3sbJQoaLt/7WrJd1HdfY5xCM/xwSAJvQBj
Etgm7n7W/8gWAVGzhXlXEBDuGNbYrLP+ml6ZIDeadg7xvqa3OJjDuEmW09BA367OOnUvRFlotv7d
Lh3bbhm8JZhyTMr4Gh4yVyinMgOw2O/NwJbLq69iGpMnKGx3JPxqZSp+ogr42qt7Rw7jY3EnPIGx
OhaQxY0E0zi9ciHDHGPJtGtxUyCvenax95uQfJu3dWSxF4R7UdcHrsWyK+F6zF+72SFYSLYJzD/W
+1Kg7KOFoIedMeHpL/iX5JD4whUyM9iHIWldppXNyw1DfgwbEy/dA6GJmdXlM8SAzO4LrlkbIOC8
a7flDJTOZ7bY/2Ayajc9FQkKvAKfyE3BrTgvkOsP4+sbkFw+FsDHrACx9DFk/cPLfZODojzbkx2G
Z7acE6Vyfg6ngbMvPD/8DQV5Uq6MpKNtdkEjFkbLdYIKD3ZHQnjJzMCX7PI8MXSqBjNHqSuYQAEv
evlC8uJmg2wOcyxEl2UcsTXWWUF1kyCsQg/R+Yp9W3bVuZx+J/dCG5mtZhCbhz/KdL9fBOV9mMws
KqzEhYTLXeQSJgG+g0Le7qdBKa53YHVhREE3PZKLcx9hJMCD3POaqL7uAKfPllUzxIUHS0B8HJe1
xxILXDG6AgyWCxR3K2YsEszZFxdV/jpau1fE5navFrDAiwZRKMgzEoNeSo7odv5756M5yTYvF8Zd
bkOGQ5CTRg+U6K5Zl5KogPF+6KK2csM3fRIVfHdxWf0zHCGy9TCIAsDHzaW7RFllEbamnHU78dnm
cVrhK+Gn6WCUuszrsiple6H6lruAB330HlKEQ8u5QoQmw3RaBFWS241/BwDcirn8AGd0gFVr1XJF
NkXVp684jkIXGnV9D5/9UX5QhR0ghx1tk5U53xCfoUYf+VqOYjKO6P3MZMzk3+n86Ts2NxPQ9jiv
7lFly76jV67+ZFakscxJKMg33vwGq2oJ7FZq9JCALA5T7Nt/EXqXnPidG20e61rzYM/Ib7iOoMXh
UqVCl0on2hGgnyM0sGtic4sLtFWY20DiczjKqt2vDH+Q2QzDOKUUtdWpekG1MFS+IvWvXRDsRjKQ
9tg3YJt5qXsS7vRCPgsAl34ZJOLEAklAjXKCUtrGfBD62ZDNv6neolNtjteskCwJVrlwa6Y0nNFO
uprP16uSYMEA90/JwP/ETvGGOUm4fayH013inyrY6n8R07TjXS6Bu/RzrxQEk24DCU4KIM6WiWYe
JlZNktSC1UXrMVa/JjT7SpDVI0VQfy5ABg2nyCw4j+0TWsS8NVtdD7ouQY0usNEcbJMwwaF/f1f+
A8ceJRhFqjQesI1mzjcwUqkOlpR0/O1QYVxHVZWFMODFXZKsv5kEngA0vYXnU0p5rRoYMveSYuLz
aXkeDmBoYy0QUiEExvcH6WukI2u58fdK0+6bJdeWUtQ/ZPz/WGvI6lgDaejTJrA09OlS05tpRUDD
oOlEvmVMdiBs+CrpXQ8senPyUdJ+JgNWBNp/TYkZufJmWYO36NOqZZbx3VVQcu1SgrCrxrfimp3z
NeGg0GN5qiEEepB7agX2hLgVePDb0/iZ9iM11Ym2slD2eKgaid6IJhrt9PwzXkRl0lQxpdvnLs3y
2AIdsLd6BuZZMOguuL5M+R4EAx7eJVpDxvduaprymW2t59OMLZedHqPXbbaSegILCEqDmWthslDz
09q35Cf/LAMlpizJE0rea4UrQLzCAijq3joBYB4Cn06baV2wOH36wPYhdrGW2TWKG3/pmbHbr+5j
CCBFl3/crg8myAxyp+0OGaYDsoN0G3XKOB4U+g2Si0+MvVusu98AuiAqnwhRdMwkn2NFEnKDv0R5
up8tm99erEgX3xpsPmFYRf6RzOT0dkGxaGKLpuqoSwkJtsd4pbvJSY32kBwwFV8YfkswZWLDILB+
K1pUjAUoiWK2cuilVXwp0b1hDX/WQ9srtrdIsBAKMVJLI1fNI+QZ6CP1XX6Fe/MTDAH+oAoXO3c7
73TDn+7bybQI8TH5qSR238BQPy5ze0BKpzgvlkDD7Zwaw65YXHxuUNF1zteK+J+3iAIonUb+9fsp
NO0stQr7gAN220uBxmNMZAek1Ch1eGE1mTBeDF8EIamVfi7WWp0UukKrKDT8v35UuK48u+5kU9qn
3OyzyXULSDQzbSDEqatS0QJwCsa7o9p37nSyLWhkN5ra/5jfgI0V5CSInkA3RlY0/iLCDODs6b8r
0QSfuZVan64UJVG/Pj5AQh5KfBEBx9I9Hdtey2Wl0Ik5uxno25ADTL4SIWPPORKiFYcidA0dB09j
p/vTJ1sBmtO3SA1kIu6JqmGFAKN/PCEZJvAXXOaegEPqtaj3TZUMLIIuAPS69IVbdbLFJrYC7hoD
Mif1sfJXkTqp4rFqPAvFP8CsasMxGLMvzilV0I05TkmyaQexcGbGGgxJ+TSzSHnAD0S/HwZBO1JO
k4jj3zg2Aw5vnWX1aow7JbmzxdZDy7hSvDSpduZgGkOelIchMoBwyNq+bQCTvzKFSvNhAdMqNaJO
zwuqkXyLjFTh/UbPN6s7EkTr4tkSEuGe53o0GoVK0jlHopDsByjWK0Hf12HQPVAIdKZSluVZaM6Z
pyQ08X2QcGVOA0R9WNmeOLFEf6TDm83b3u2g6YmyCD1gZC7Zc0mrVE3K8dwV24eaFARXaT4RRrJ+
/thIrJRXIGzBkgcegQ3aQhqEhjphiBZYxSaAPQWG/WGpAl6pzUrLVshXgddmpbq1vrzmok9aZJyE
ejxTXh8o/dIMseLsQ9vyMZl5w5KIOo1gtDemgu7ywjdINXZ3cMWHiyxIxQ4a6xtqdCX+wt/aoo6B
nwCQjpdzOA9HVloRJL5OEU+GlhrVl1niv5G7sNN6w/3HvKnXVNYawNT3CmdKIAFWvS+789zwFUis
xfmvAuxnbCFYWgJkWwf9Zn08vy8kSqSftAj5DvDFIE+IRqZ+WZS6HL1vu+RdKV4k6nXq8qO8jort
F2+5AawfSlEQMZuZY6+vzjkGoH+V2loTthh7tqWe+SNsosACU7vrkPh1AlBUSAkZtR1qlLyuBBrQ
Pca5OShn2vUEPAk2jzqAQoS23OzFCx1Luyv1zzM5hbAHINuU2FmTH5GASklK1wV2kU0a6rQp3Alw
tXUQCcTrDhGOZozWWuIG0mkMKPIo8lgJI5Ks7kjxnHtzfm2WvHapk4gWY1cATL+9UFBljG7RHY0i
A+ofnRMYlpeaEzpsre/Vo7JS/Za0TpfRMdPQ4XXQsjtsjWBa7eepcVFDzalTnRPadXEbJSkq1Zor
V1U4fASE3WJQTJp8UplTbRcTx6useSrKjq3K9oepboGdO650hDntBTvdRH88AI1FDzSPrm06zBUQ
OGj7TqXJhSLoGrsDyrfPjx7xq+tXTgJiyfFZvIv9auoEDu3ViTftA6Wvv7im8K4Xc0+yJ/aQ1Pbc
oPA8McPN9ZawyLjsYAT+qLpk7kOyJKBW+NoNXOV2GzlIvU1Ohlpjfqvh8DFnWW8J/tWi9/BPaiaJ
aZegVyvbeOUvsAPxpCvABpgA3CdEHlTvVnnUL/lj9vCeWnHRc+ceF7yqoPKtmaeFAbsBBKmemSTz
L1805BgEazTvfP12/q+6nLkNBCBoam60vN4OjrpjMLHV9rPVmEzqDiZF+e8ItzIbycWw6RyPvh7x
ro2oejgK60QqL+0+LZfUbQkYDjAmVrOSJwhLwElGhhYHR1084pgy7VDNgGEuD8mJgBot2ZMBxzvg
8bUca6rJNVFMVP34616mVKVOOVjdE2+armzdyPEXbUodWT2S+nRo9kFRw5CPuK9IXUjlx1VS1oLn
nmhQFUV4I8QJYEj7ZuHHFvSH4U0boAQDfBh5sr/5ZZcybDdU5TfQZhp4Ne8hnnFiymeOZ+Mkj57f
umNfdB3wilBgBR0EdqgbujAW0gwRUJNGSO1R/FJwooknV6gIhG7uAv3JXO8ImrWu85cIizW9r9vX
TJlfckQzMkuv3r0Sn7WbwrEybFcIX5flji7qMqmylRlwOIxw6lxxoH7g4zZ1HgxZzfPHLrdi3FIg
OU/c8a22CdiyKAMH2aM+I76n8O/zjh1ayipD7bhfTHrMo1NHTEyXdc7ohngcLjKysu/g6KsqBxGu
BSrl9cUhoLnUKj5efQH9S31tIH+GgPgHnZ4WAoMVPJsSnr1SJoc68lMwIeA052UQP2Cnyq5zftA1
VG3cHxfk6i46L8hPGr9pO0jvKNb3xyfJuox+CSfh1tQSizTX3Z1xg1xvkkXQP4XnqQvM6SKL8M7R
6eLPp7AE1+mlIX5fXa54DyWjAEx7OywES6WTlmQVzkQz4vOcgCmdjwlTHbLtLk9Uj9ksDEKKCcrG
ENp+lZvPK3Os9A9AF7PtD1R3xpgrUlTGMrvMM3Xjyg7OlXma/qK90ypQU1eJIPJp7GWBFgaXa8VY
xcD0JqUvaomtVyZXcWnkIOVBx24cmm/1BLSFJSMRXnpsouIrsTpzbiYR+3t4MDcsp3JDlOWhQiZN
oqqGqxn1YdDTwRjWATcUNFxWHWkk0fVIe7O9lhp3XvbkR2bXIQXfXCKdruZHkMBRo4UPdbzh2dhE
TpM0pPJ72POmuB1KisWJhQGeYKOu9FRNUX1KFKX/C7AdbEYVq7tmr7r3y3dPckTOucYrRW5OPASI
v06YBebucSauMNq1/PgDefTjYJ5dcg5FIn84p8ksoWFKryKJc/d25IPhlqRV/uEoEwui7agBTDKJ
OtqgTbL0ZEiyIuYeYUwVDJEcpbWQfcJ8MfvWr0OkIGW1vHh+It++fZ61uqoMLlCe3PW3+PDEmcgJ
FjCpwfoxz1AMnglv61+phAnHpvAPJBUTOqEoKrwIWy36a78h9VUsvqtL2fKjq6/BNLbzQF9IuQ36
n3o/aIEymZnGPO0aQFqkEGfV6AJREZRCEiO6XjAyZE12ymtus8zMQ35WX9Kpy61zQTiExJy9Xwdd
xYxZcn7knSBhSond0fyLLDsgrFqWQorFhoa4gjHuh1ZYxypjFu8bRW9CKc3kV3rmsyIUeBIEK7L1
QHIc7MFtqGkt6XsFp9O/uhNZHIRjYSHhUr1olpH25ahUZ3xmonB2ur7xnMTagJajt4uQeUMVq2vn
fVYNhaUf/PZOkoBwqBxYrXaqYehocLn2lwnZlf+GIQcCJV9fLKPex2vf9VPMuqxHairjaJUlexA4
fUlorNmRLtcN123TINnUJTPSAk5ZiByCn7grHCG60DEwE0QmiBbUf9DPqxaWdu4Bx9qvUxo3r55m
GbTWV+phKU9V0/iaGhcOwl59WSnN41aKYT7ziurxu3n6vX69tXmZNjzKQAXG7oHhElhX1Oe+pPR0
aqRd80cqOT3P5rjo0v8uJhmwFYfsIj3wHD+NbXL/5hKZNEarQoEK/hBVeBBqPxyxUBsrUf1mjr6p
1+62ar0LJ7ub7qOc165Sh897i49euknfM/kpmfmm0h26oz7jTh5z505ICTkpqP7Cs0TE+3IIcsQZ
osq7byrZd5gaxmdPB38Ulz0oBIhrHSCJ7SQ3R1j3+Q/F2ILsDIdo3v4ISoRopTCIUsM43ga1XH6I
afXKsgWjz9A8gL+WtM4d5Kx0KG40VtzypeQ8FQnEgIvN4iBSZfx0JtxtOnGWanN5fSw3qYCfv/k9
IhtDro6/8YL7Ud7oPqCjMkXOgfeHCoTtS4tNcgfs3qhdnXV+EiqJJ15qOpn9St3tXYw69sQvOwhX
+AmE//jnHn+hz7Al6k+zK+mPpou1lwiBcql6tLtBFBa5Nxj1EIE1wo26jujRwXNBZMxbzoiKK5hx
1I7l3NrFltN5wE150V3JJHTQAQYcAAl8O7fv2x7WLnvleTiflDduBDNjf1Hggqd7GDEo2YyeOQRS
Psaq6KdEvxglDSYgyDN2Gv7mBPK42IEQ7b1oZsHOWOhASSjGmwnu2eEt4PiRVzWXP83S1E19oR77
Le7wCht9tO4QPiTS+AsuslYUAhW9Ribt0XvfJGs5g6ZIoRqOMD9+EsNgldWBwDGBFP8DXAtSanb9
o/ojxAZUTXIoY9kyTfTyod7RfrtuhpYgCPLaDdjErEg5es7PeXTB6ie3t8VRe/zDptZNAiG8wWEn
BPS0H8YM7tifszADGI4YXBbAMiqI1kqp3cdyzTdDrQ7SRGSWGC1wnFFRKqpc4aOo1R1smKrRg0KT
1JICnuWIo558jDeOcrUWJ6pt5XF65oaBs7P46XUb+X2v0S9zA7BCnI0Pp1aC0qpPGzVhiiVu1FAu
u3cuHyAmUfHKlu/maBkGgvXsHZuvfAlpUEWY7hoClRmUd9JYC98Ti83PF8YLx0s2VYC006MMbcNZ
461WonleNelXlr9OCZdYDk+Wjvao+Yiv/muJIJgDF6hghp3JAEEQI1lL13cazi9djLLjGsfmZUu2
C2j1rhMSoknminh71rtARpg4T+nMz1oYzM/bsuJ6HSPdPTuaP4dGh6wqEpDNsin/L+DSQCU9z2AW
PzM+hZGszXT4he4KnAOnRKGPupHGILDlLOT/8/69eJZJk8P26X403LCPiC473kW62Kdy2TKdpVyj
yE/lQKcy3IvoL2aBVGq0YrkHBhP/K6i1i1UuVykmlNrXHnDdVBLYNO4PeaKM8nmrljzGBD8f9pZa
D5FhcdR1Z6CebEu7a3dwlzNrTeBrpfeNFlPru4Kpv2c61GOWeoil8rJuDejlebBTJylYPcdgq6cF
PrDUUCaTzpM533hSTDcEhIW3HdOIgQ5nuHeHsmZrTuWAzOL92Kg+Xtva1Avb+FkgABQTtqEoY4T7
V0U9XF6yriHSm/sTJdNXqKaJPbNJobobeBic/UP6DYf+GFlNdGOYJCGacGu8Me65iXPu0Om/6vuq
ghU/mPvRqa4u9sMgTP0S8Tqhf3Fd2k9VEcmbABBUCGyNClfM43Ft3dZQjXl8x934oJQc3I2BWg3t
J+yIZzYNBmqMyxZN/HOWNeY2y0IFN18q0P6TQKoJOtSwnQ1CegfTpdlKpbu1ByeZQFs9EaVfZk/J
lpygRhRn3yPn0fdAQe1iXW/Ct6e/bZi4KyRfYCo2zdjjTAvCwkeEWOU5o2AhyOGFdCirXQ3Xea8I
IBaFe+lZYgNIa2YblA+D35Ei/Sb7fxG/asoCfXraMcPPiSy7SHXZLhbra0XNlOIZUsEjAJdndBxT
28nTi+mDYTB0PcX2D5pokdlbUvRSg+q9aQI7wbC/6mzwTmYU65uUvCZjm62lIhCGZ+tOvXktlk9t
rl1lX3u4MHCMuYmg1uByJZZgatvgyfiOpqjMGwKtJbWsd0BhPJSgGuPpOOQUsClZfD0yFxIWG/3Y
QE16pbhxVvM8aJTgT764nZiLst7G4AM8B5OVTRL/vOhFcMFT8+9fpfPp40I57xJKj+a3Hs44794O
N5ivWnAUbiNsr6Sdoi6qjxK4hKW9Ao+g91ar+8vcaXUW4YFNEZwAi73+3XNI3S9CDhVTKL+6/U3D
Qu8PifM2byfwpsPNGfNdeHAO5LfWXALtNX2WT34g+wcpO1WiZnqlkxjkRCSvOlxflpPZ3GAUosnt
akZkbZ9sDPdWWANq7C7gsfeKQsM62/mR7lQVclaf54d3WTFqNNLWaOTT91OAkgJPQz5k115Jg2W0
5yb4hNM1sWuyl1It4Q2i3fTtBo4dgaWglCweGuRzBomaRmpNB890o7+1AxLTERCUSJO5xib+YBfV
liK2dI6PE8Sl0yJn9sGZF4xTX7KEUAhLuw4zodiuvLdg2rP2iwKBmCZk2nbMxEm4alpAdIjeZkK7
6S3hE4EvS/n3N8SV8aSO+UeEpxzauisFvCmZOlAbvP0stuo5TpefWdxDM37Xgt2XB0sYhgQzm8KH
QAYew/XLBJG+yC+V7M0/Ey9RcCC3E8boXFDviCk/Ct0g1F9B2F+wTrcf3DuNbPgwg4gQh8fvfiDX
snYh9TpRdjWZbOA8oDTYV/1MIHiTeM1R3YoQ5OlK6hYkAiILj7V9QXOx78ly8y1AXUR+f+wTotAl
d37uIezVqyZsGF+E7sdn0fB5w5Qgk3Pe328ab1jh1kEfLYtwPf20dHEGH4DFp8LDXpTNt4SQz+hK
9glRY3wQu+UaOIVFgnO/7h68x4efTLG19o5lf/ZXV2X4GXiQ6KZVPi/SAFKoZ+86kqmRXR7z5LOV
WeqDCM/T4kIwIqBSjjKq3lOnhDdbDZ8Um3YE8vE7m/LV55EgguSUz3ZQykufrZMaghwNU1H9YqJ5
Yb72eUyFYXKTLu1S1KT+oBRhX+mN5t/v4oQgK3nxgc//sZADLqs/Dn5CI6baDzk1qGvv8YsmiKuz
WsIFPVk2/d2ScXn6HQJLy+FSx03q44LNcc04nYwsPflcqljgsQhoLHNVaGRcij7mmsRtlVIgo0sJ
V//o9YAnt8ZL8WpLavzUqR9wJvZUUtuv4tZRBEm+t6dnzAsgr3/UP6ljcUGF3wgPzsM23IZNG00b
6QhuS8mm8XFWQxfrRd7sB6fCXez2LM5jr0LEQPSYgROmXQMXvNg5EBvS9uGqg3gjbDZXHwessr1E
O/avCaLAvZ5CxDNsAeQ8qnlpvfhhMdtelaFKZRQSOQGZn9HDhuzUyB50bOAXdhc9QY0gWlnyISN+
P71X0uNOZLTNWMF7q9AvHaCBuQn3ByXE3VX6f0e53CI5rN2HPNAvm2qBk8qc2xAiNDGCuFWMqJVu
5ylZV+5jWKJQNjDMnpoz/2qGOez/ZpQZSUQbnbzYGcbmETZI1UBZa+SNxm49jOIeSDcLQEsgMGJp
8Zjw5ZtKV3tx0j6ul+QBJGQSCAa/hilWSTsh+lvBNHC5x/VE/YG8ZBLkpgCZB6alfJTpJK5tSoWM
48BsxN6N9+Zd6TfQP3pFVptDp7oci65vgpQb8jqU5hAEwZKEWxMTHT8PuBE2pgpuaAO4nO1jmo90
Ku50QXooJd28qzWCVbRnVvDn0PlsVCLrAE/hvjPCG0pcBiIoy37x2vXrZ28seCj3JCXJS8KCUZKh
LmRAnQcwFxMYe2HRfeKzDmz1CuRbLtLuxLxJXijq/mYYGu4n2FVV5awFKlE1+yON1cXqPQttKHsP
39qxxMRMVQQegC0lvSDb4i1zKdW9nYTfEOD/F491sct9nRnGW+mQrnqewTzvSzWrPvM/T/+FMcLE
whd79d1AEivlyIZ7gqDTAwfVWGkh1m2yulTQhJgsOtK5JbyJps7IwZA0sZDX1WF2Lp85McbbCLOz
BZwzUZ5/esmgdTJSoPdt5Cc4Yfux33zSPaf+HMMmVfVCj5dGdxIJF9rEPcP+lTO0ed6JkXX3XE7K
hpIXjmzxT1/betwZC0MwGWlJC1e+wvJs2PxO0wjPTl+mfkyZh0jzXIkJ7g4Cu48wo19VlREShNPH
nswWXdI4JL2QnAgSI0arLE8ZAU7Cdz7eWVsqYO2uwu88dbmI46Eron2WNso4TDS494Kvez6GCJ6d
8EKAmj40yHhNjOFT8mlKhEly2qoueb4Qirk+9QboFt/ZvLaQWb6/wmFFE/b5puDcM+sdCiJLcJ4y
7xY5KrjnO1dGa1uoRlEQcWjc9QaUqmqtsLtlWSioUvEO5wYT7Qzqf3BLbTfUTOjWb8XjLdFWsNlX
PbV37cWyjOPQ9AE6xY/C9fux5L9BV6ppInr2lopjJdlOcEBtTaj6LbwO4SRGqNeA5Z431fLihJdA
et5Ro0FxATDDGK8aRwOM1fH2G6eFY5jBs8KGgTMZbyj6xANsLOyMzdqDfrrNpj56YyK576sYz0uu
9doJDpMuLHsKtyVB5q/8VQUoOXkKOSquAi8d28uAP7pk/66wgZEgQqJd/9NGLlXutKLcJV2d1A14
9Nc8qxUjaZrTlJjwJ2cq8PvDbGo+HzKfDI86YRQv6VRt3S+f63LWvaA3BrSkToQs0opFqY3qFY7V
nlhnFEsrmAHcL5KW9Le79e9O8guU9xNuCkEf9rwIiJbfMgJSywlkzxldsSHEcxw2xJi+TjWhT50g
PS7GnmMFLnLuDhv6yXGyRPmN57bqkivlhsSvcrISdjEwLuGVRxiKbzmMCAxRPMFnzTVDEzLfbl9+
xoAQ7RtGFNVHEdh15O4eiBhnZVaU/6gJmyjFCNcoHdxMHTs0XiOnUI0Kl4NI0axd4BdfaBIyijn/
LCpW/YFT3ijMMOLxxiklX9ZkRzXm+JKtqIFOLs2mI4VmFj9nIO9u2/mA3/LF3JqDkLv+PhjGKePg
xFg1+SXp+jR2vnOFKxAAiI4YTmG9qL33H938VKks3kAdJj4+Z1Rwcwo7tShsMIrFzDNfdl2HNcu2
wDQO/RfIVMSXnm/+3dpBEHqcb5QuCEtYZn1oJT4tYUO1GzxbM+8/s5qYoz4c4bZxAONj3/sz7bSc
a/OU+248UigFLyb2kIqHRYkCyqq8W73k75gQwhOe46kQIZm9SKewURmo3NMJO5qv2/SM7tF1FlOD
xLfaj/BaVTYanIU6mFT0g+fJHsWRioK+lAuckkNLThmMsFejC3wtvBU/fD2rAtHaZZA/oZ/rOBy2
6c5ZuOaC+6xZe0wuQH2CoP6SGc4FNxcUyxpo2gVCxD/aO5BEygyI51ycGsyts5Ye5/A+4s1hgJ8U
QwMs17D2JCt/Yyr5UziYcvRRY1kR6k8czzXSCu+aRFxtOTNCDUR4aLYqFSzwAxRKhqapMbFW5dLG
UIgDZBRca5KH8y998u2qIbtal6Twu+yvD7GBIaa79xUAoEPRgte0omC03UxyezbHsUMssMv2swJ1
tYDkl1bR083ORDrYjwcEaIZhSp9pXZp0WZ5XtZ8ID+i9AdIVjg1r2iR+KVIf35JmnyLRZV3AXnwu
ZeoGwIveVsOqBJeh0PQblgGfAmEVCp/7TrapZfNdpY+n0N0jOb2UwKgGtr+QDiFTSXPK9q88ZAut
tjD/RuVB1Hx08Ozx0UZkhBV82cI1IUQHlXiE3KID6edAaawOJzGpPQf3TixIrpWb5Vv6wIPgJQIe
CdH/3pF1W7TyNl6tGnFpGRmvwM4wcP88elZnJH1dLYF17Vc1jsoseFxQDaQspUiabDT8VTqo12mI
c9Y8jv+FoSn8+wAwaVq5ly4T1hNCcMdBnMXi6CFfQN+9c8ePcTJSlAKP9C3hZuYcv+7lA9xvemsN
eppbSaqOpjF9L6WUvUu8y1fgzxBKMovNw1IoJ70YZ2fGUzjWE/5T6HASHPKsIZhQ1IF3z4l2uA12
5CQSiHkB0pAzM7yNuILvhimKsNTZ3J01cTDJNwTxeSptBrZfLp6pT1xzMBjZpEU1/7NfPlZ0oO8x
XN70pL3YgeVs31X3+17NfNKDOZ9fkpKlqFTxNX5ySmB9UxDoIBl9H4zsDJhV+y9ZkhjxIjNxzbx8
HnDnurRrsT0hIo041SplccuwVPiCgeT7PHLtHCWOO/w5Yl7jpcnNsvNc0I1vsPZwL1rk7AifVqn9
c8UI77enFvUtEzkRPwjar5E9a3etm8x4/YxazTzacItnNtdwvdlVt2m3kM9fj8BWaZCrOBCefcaK
iKQqDxj4wFYUDVOQRs+8pXSxUsy/hDHjs1RCEk5lEAgAk/ba+jpOvgmOPUpiEJzpjCKcNkKmhroO
8qQuS2uYAMn/br0zSl06Nf/xS0dDSZnGPjqAjhG3MIka/dH9Cv0vDbQtf84Yuzlrk2W/5ufarAXg
C1odv9vW/Q0Cutdy+Wplv48L55B7+FBVZZw31YowlDJSH+Ga2CgGaeVoNerq9axyKYGZcF01Fbmm
rUX64typVkgpixpf0dbN79mZGy9mDPKJIL0MQ7Bv4IcR1tgtKY8bQG5kU3gu+NqqekI4jGQtpru6
/XIDKAVeGbSnlmZ2QIybcn3Tos5B7WyVXlUajNM44fn1MVBXjoIicU3s1E34rtHIJ/rpO8YvG8bg
X8Ky3cKAWXHVK9Nzim28rw7haeasewB4M52VOXiCHljKQgNv4UNXzSbxawYArySUPjUTSrWOUlSZ
jwgBxFsSfwaz3bMg9cmCRM47yYR6aAWTDF3hY/0RelTv2aTB59ysJHICyxFbD68kzceCoEH6iYLF
WnTFb4htUfR+51unROb0Yq4ULyQroW27zWKVngDy3ERIcnFyCp+i6hVNVieEB4vDXbcarAzlO0Mz
tu/LZ14HYqRpkleFO23DSaja4hVwVtX+duyr2XV4diCW1TWk7Vab8lRbuI6XKIibqdT4T9XUG1C7
ge6JZPcpsIGoZnOYgkv/sR09Z0JZewDyDvlkTSelLTK3Eju3c/Ej+uKBF9fjWNm+kfZvHG3trk7O
G7CROb1zg0BLmm85yYdgkB6ZiRWlbZnBIWDKmBV2o5i+9E+cDi5dUODOD8ifnmOs/5XWYbgqrPH7
5BmI79Lom+wLsuls7ng0yusKdF0uM3hNkT1M3NFmwppqKr75nLglGccy9T2gfBW8yaPpt8n5pyqW
dELsAxxG94ChCeeXLrx0FuxyeLlhNvBBP8xvdljNs7zhhcCFZN0GGgCoYkbwtPs5B8R8PIWxe8C0
CVLAayF7bsLoHJl+mZvF52juCrJmI0SeKFXTO5OqoLmk+NnTEn7kF54VU8NJ8rqnAkc4nx+Hgf65
Ktxgpze0kDOrdum5J1oZiOWd4xNZNcRdUEx3EpERcr16qZCzol9M8STtaJLzD21H3+vge6VWKyLG
4L5hJSxuohAGbplZte4P1IzlsJW5uuZjTeM1aq3FcTyl48IiFmSGG9IsaVhHjYVZGPJ+y1HEj4KL
I0B4mIsyGFjsaQFBsAkzus9RnqkUw1JFYsThLftlHAwyq3A6r7bKBr8TohgEjQtJgLfBeK3uzUTD
9bqbww+OgtW7gzZznMd3oZScgS8+SVqX6GAKiPOx33EAZD5sln/43/gMhf36h9lKqPZvUM7i+ZWq
FnY5IT5RXgY36ELYksLtBjcubYWd4Mn9pXg8G1/A8V9wkP0X4mP07GraVnbjjtiN8U/8uQtEzcEL
NagyMFZGav23QrZevkWj7R2NGbEnrsNHQFLEIQLFJRUmJSfBX9yC/j01Yj03zORfVCHqsW7LPTN3
HiPpuff3rpg0/EbVpv8VOD4tJBElPXsnw/goy0paq5sUz3q21c0uMHYYfcsCgFxrIwDOeQCEgp9X
fkjhMG948armul7zaiGhl9Si7q0fzbeqCubZworAXmFmUIjPxWk2HNXVEYgOe2Cb3cf3gCP7KQ0C
XLTUkcdXiKTk7BtvMlhYsqZNMlmamv6+7plx426DIwizVG0DVmyjtWmN52JRomKqHV88PJK5+1hc
B0L17WYhO4+JdqZ27K3+KW4WUjMNinRDRxaZOfcoJMYB42s6FcnJR3T4uPCmVomodizDYZtk6kIF
ysWmtsRI71Kz3J6TK1gLHq/qAk0mi+dBE1kH8gi24QsfiDbyo56iljWwIPChioFVVPER2dRPYvUg
j4vpL2lfQBY3G/VZmRhyN/jP54aAKrU3qcLWHS4wji2R07IdiwSvw5iv6GgTgvQw+nOyVD3+hcis
g3BYpg7MxXM87zldYz8ijPO81Gxl88VEgTKuK6BVJORwS4nHj8Y/6/YKq0g/IdTtOoMrAcnsAOm4
poo6vjJjwmoCLUsU6+jTCuOhYlBJHmKCEZ6zkFKzakQRcI0KQhmBRxNdHAoT6TkWbSGDDBDZZV5p
7a0u06YvXLcXfP8LzYybTaFtkyYZjqSE0eYQeNyFNMFK7To3SZMCKoQxPBhaav6tLEHZDo13ijsO
CNCBZNmHbGCaWpX0plLy8Ipjskd3kMc1c3QbQeUKUyKQXrh8S2kau96MTCjjfpIPSYAaY8jsU7Nu
8YocHkaT7wj8m44mHkgfHjSISzg0N5wGwLf7ybPPyv/XZme1w7dh+ilOeMZuEKcqN9kuhxeLeQM0
ESeJJ1wTlQyuCQyQkpP3OJe2sHBZJi26Yr3ZN3jmVViGnRTC9Qe52S391C2wauHPbJQg4FPKZMHy
9rHZ8PJ8x5B473Iu0XkkV25VXIZnBNVxwVTWOfK5m+ecqjOSGgbbyCWhIgVAUsUmgKN5SpmKfC1u
0HsPysgyUsw1tx7779OWCvdAipu5/YnvahZEN0Y6Ihv2E6Eyl2IoZ3vFWqLVO9s9Jrx58LmTLq1N
YMrGmjFTO3T3BKJTJ8D3yvrgRBzFHgYyzXZ1jdnR/BiccRUYb+j/dA0KmPoFSWY1LWUGDkIV/Bcw
vUVOI/05lyUYOo9Ngvb4MVguPpIL4/UGus21650qX6+RUSjhcpbDq7c+dX1xWflcxFha4s3ulTGC
FmgzSdzxokmjo7TwHpt2oxxlE4y3WPAAKhhPS9pxsQY5bs0PebCWftOnB1boUW46w4T1ERNuEQJO
BiY/ugYqPGt88CMRTAYGe99/E2eSyLvPBChzyDiFp1G5T3tIx+ml6Ow0Uh2lXDQ1vDVOtlg7SYqj
fTV5R+iz+WiwJsNsbu4wBrXkYTt94crLee5FdbyMfRL+Y3uC6xLwbEEi6QS2IZrK2/Q2P3yaXy+p
wgoXJpyHJpY3KeISApP9PAA7d7sj1SCkTnmzfOo2gKaoIQPYxSY/EO/CxZSHie4NvhdEEv07TEro
QeNbsaz5Adno0IhwMnm4ehuxF3sYQYgMLl5o3lmP7r0gJGd06E2d6Za2JmqXmJS317aWMNFDBsCl
1mqvXbYwrwJw+mxEL0Siv0ysRFBE7MG9gsRk4+6KUbk9Hz69KMH4k0+4YvQZEceZvsGwCOcFRHkw
9TgvI6B8Wo+TlHRIF45t/YxWixP5wHsme7SDEyPvxrAS+QlmlzZqRtKOTzPwVjwZfTCh+XI2l8OB
kc62NwB6cQ4+pFpq2N88gR6HF1bVCyg+gaiB0HWqWOX89Qh5Utu9S6cSx83y4jNHoaWq/yoHE7uX
TPXDuJTUqskxm1jWq11VL0VFUCDY+zbshj6JtEqkgMnnhS+OXVovKqvtXXWLk9pNorHkn7hAbzoC
NQVDMbZ1q9VZ0BTPUGESD188TV63Im+pPJkCGE+3qz0Aism6fj97Q2jTgholJ1/Gj+ZG7UtuDxpX
TnXuJ0qIIMGlZfl1eFXq6WIviZkZXzzLKuQ7eTq6aOyXTs5wtKkLVZABFo2yoqY3L2+2ifGsVQDJ
3OvF9Bphvz6X0Keq7EtWyN0fWzFumrSZrzf9xABDCXa5B4nVmCce0abv8CbFP/0Zp2N0OufnoB5D
zZbEg+KSYUFNLqduBdZDz7ueesbHxjAsc2jKTrQPECY9iCaRO/bqz3yTc3AGaBFz6fVChhD3LddP
OE9EICk+pKGKwqVZuOQ21Kw/RKyr3E8KZc5AASTdvDpQW///1/T/FA08+4kjaubuBDAvPu1X9vzI
sF7qyc9n+SQ7SgGpJSJNYpZ7kYRETHFix1wN4oovesPiQOo4I0GN388ktGTK2+GS2wdH1/5dl5CY
/tUtGUtVefJRdhMbJTcAph0UlSjBWi0Hp+dtFlo98lgenQuOkeHimR6KC5a9W5F6wdm7CMrSmxai
fu6JJrTvGATRaEraHWm9/8lk0ABhivJQacWhEcwJP48TeCRwt2fNTZggswJ4GErzRV1JSYzFepRw
uJRNNPBBSffOYhQ2MEee5jbILLNFHmgMbdFlXJeTb7ztVA7XLmncYYqNQNDOtP0oyAJfS2J3iGD6
9qv+FeVuBm9k/AMNBKF+jxKxjLTUBH7gc+UDoIHiPAB/n3YRIxOogls8c0CKSfq8lkrns9AvHR7A
pMn7UNNnxPssvXASCULFjBj6U8ksZGV5ZxtnrkcFqxRZxqf/m1ANdGIrRHEYnLeI2SESrAuG4/rs
tqVlyh99z30qLFwrnhV8FGRwAwXjJoxp0ThCUf/XyvCIShIJ4VesJy5oQ+39mWgfeg2vP/x67ra+
Whmb6sUBd0/M0uYRYAzg2Qft4Tw8IMpclVvjFwm5v5yB0gVI9CgK5gNefvPlLkkXxCq7aAHPeBP+
zdwRlgJ7G+yLqCr8M4gtciUOHu4vUWS/NFUyyZ724MSMBtcS4B8FYEv6LMUBqZgH45geRGShq+28
pNbJizuvUrffbK0dUK3a/ePp9ae/osVNNeImTZudlbsWaOV6ahbG2SgZYei+jbxahwPqQ1qRmw/1
LW2+cUVrSNYkHPlJqr8zozZzuT/6GbgIUG0b9VEIGdGEDiJ+qgYLMYrFqMkOglLnuOzFXbM61mSu
TY6hV2lB1l1q/FunTvE17BA4AzLnUsDmcP0ejMw4AUJQqEMjz/Arf2vDWTs7lbQIqUF3p1wnNNK3
QUbrn5EPkmoCMc/jgT6/EISJH5tYC7KGzF40wPhO9j3iPdbP4IzXk2HPnUZxEDVCi3oGU1gsExJ6
cgUkOSvAmXqu6fy/DGlBXlP8iFO8YHpEbbtKWAKHfkutJM2Glvlkz0wQ9V13k95igHJ5/ZV+Qlwz
fw4g3WmTaURFMcsznhvOjAKVsjXPVDYXpR4QVTQnmTPeo1eH7aNskOKCIYjn5+D6idfug3GoDoHQ
CfsIe9VxFNrQDYgPFglpnAhq27aplAEnQsQoqvhzZ3rj9Z9vk2dWhLPBd6htBOuHk2/pR8vOEGsN
uj3bPI0rySMU4PUha9iCMJJrp9Te49WtG47t9u4dgzHcGm2C0gW5Q8xDMDM2QaRIHSQisDT3OxUZ
Sk0x8xv5xVXF9wI8GvjXgR7hwTN5yf6iPsd2WP/JwVClV/XIESozaOHspFw1Kr/goN8nAmUAvx/D
18rLAgAbrHdFHqC/QJ7fHiQ6EnWDmubJra4DUEX9ox3WELHm+w3YZuztvZAw1i7Sp3br7CLShe79
FiD/d3asq4UeswkmIlWTQ9VGoqwdBXq5w/U+cEbMyTrzdIpYc2Z3hz/CT7v0gteJnhWlKzm0tiDm
aisVwm6YqNcnLF4KmcFacwpdx7RwfJ99mU9X06g6q8dcQt00eJ4irqSjUFOFJfc95tj+ezF7/YDN
tqMR3RFjHEVAvx2nVvwx4Vu10jFgOOpFmGN1t+R5mI2I6VHhaxWbliF1lSWk39xLeskx2jo/7hDx
JVgIsGnQH9qb2cSiTPGVu3ax4Z3blyr4nA7NiaXdp3Ylr42dkR4m4OG0RJIaUlA7amtAXDR3+HCS
F3wbOUHIWo0Q7rsRgU0HwOsCNcqzs/jUfomC2xajP1eMsZ2dP7t/JMHgZryOGbjZbabZUIKvPXn+
S9ouElxwv03C9RxOdyDvHHWZVOg0dHmbeRvo8tIlbearY8MLPUsznRl5RnKcc4WpONv4V4AnoCS/
icNO8hyxNLErQ546CPjdhoiBYfA9ixo/O8tf8qNOEsZw3PMG0o4z61EZCS5O6QsQo8H5TZv70RUR
tI/wpkxxpkxyIr1w59V77U7EQrgoe43PmECckhRsl+Tpiot+JrHGeAdUwQTRjg6o+B5GCi5wGy97
C/TIfq3NEEBxpRSxisuKLJftxrHX6ozNWpTaWfeALbp5lTkidzgGkNG3dPLbda9y5oO0OaGkQ3he
Z5vlbl0aED0MYrWgNg52gKMtpQquExHZ516z/A9mlXlzMwYNQWzvSciPAws0x4gwIEdyC78XtbI8
xvqXeCP/UsmDWmTgN+E/ws34xRZMNkYLNp/pow+s9nY74C2+5pVjYsWg6YypaCpmygwxhEHWxKWv
AheJjFBqq3IlFkV5RrVtdjXNuKMbYhSjK7IHf72r52ro7y7Ti706Q8CPDj6/zBmza3dsG50/gk4N
I5FXmU2rFj1uE/7iVxZUwFfPCnrGg9Ch3fo9vTxVeO0XmJle7jmYiGLl6jxlB7isWoda7JD+iOnO
uXCwpXowbtdKlGRpH0BHdJbHwZGc0+mXJx3r8ikNTvtdXcoEImfO5zqv0iFdXYo9fRhCzr0TqWcw
5/j/IgbpQCBUz0fiYACi6eiyahgRgTsatc/F324WeOBVPbPYZqobC7+2mfxnpX+VdbcQN4v2PoO7
ORXjMEq8wa8P1YAdDqgy38HJ++fen5kfJm7HDIMgirezU6hJn6aFiBZlyOxM87hdT1IsQeiw09Ps
fzerofCdmawCBt2inx0FUFGLI6c6PhS6bvZPb5yhF/Dd1Tzp1o1AHMciy/QL1QcnI49OMN0ccY9f
TE10+nw9/46D1Fc2trFyWSbR/wlguhbWiOi+8oMj22y5p0iw2PcrzTkTSWqjATd6rOgb/Ge7kFb1
YoHHFZ76n/bsldgfvEQ1i5aGVvweF+GThL2aXFtK8UBS6Tw6IpX0NK7+X1npZDXT/pqh7rSFVBfA
F+qk0pqQYRxhaeDHp8wvQ/0OmP9YSKJC30dg7fkdKhEakjH+ViJYlY6Obvxzjp/+MCBe+ZcOUb2k
jT0oKWQXLSZYfqtgDd8T5WKexU7/OTvPzYZXAtG4WNcC/V/PNA2O6xYDLS4mEiBmxpNOHeyrwpXC
yf66RyuZHnU8a7yTgN+Y3lYKMfWKMIAL+Rnew1SBiVQ+TjF4h50U2GvWxvSTUJa81ouI9wuklRXy
grEdUmWB0Ur5AU072/+EHYbhGaeZKNxxEGyyIQx2IlEPdo/xsgzeoZLN2vdUI4t+rCqd4D7VWP7v
+XV8b7rq4eUmo60lSP3H+nD7bpq9bv1UYWc1G7Yl+3SgtUYOLx2T09FyaIQWybIgWSMf3zIqkQYy
YuxeR0DrU11D6cT0M5hBBdcwAy5j0XAlUZ8F3TJXEnE7epc33lUsHkTTg16igIe6+DO2wYxXjSQH
He2eSD5sCPM/Nt70CxMYaFwp8pRZ42/2m6p5bEf1yYi45obq2sq6roeLE+RrJFRqsVbqW6D0OswJ
xNLeNRyVjN91ql7kT1Osmnd7aR7fhoWrmWsnoK0hmH8CbwVnn1HuBB83KxCJOIbLsLZDPPNmnOsh
Rhl/R/3k/HFLtBCRwNzlhWPt4h/zP5nueZrZK/OWOt6B4UBJ1yYx2XR0wiLqbkkFjtKQToqjaaNV
0HbjNAfB7/fWmRxXo1b0jBctGCjAfSmnmlohu7jnT2mTQk923U14MqDCWrfrFFaBgMM4yNeNvGdd
TUSnhsPZOnYhzPXOBMK1MDbZZf6ZVGqE2be/Ju4m/ij9nVlcgr/yi878SSdZ4yBFsfZOkBLkj76c
M13JftRd3U6oITclVX8qBvB8Qn/IMAlxgVOmnZZjzcxBfWhze6fQ5hD/rMI0TrIND7VChnWk40/X
o8UiCmiFCEOmPquyDXabuwtX2NTvESL/ZwUxZs+7hWNpTGify5caFd7QTai+wLwO9VnoAixnaZ1g
9ufLGBsb/jgrzr+R91tQq7knatSntKqcbgNooI2BfQpPCncfazriVMEJ7RmIF8jfzIhLxQ8gaJF2
d4lLlY/NrrL0zPy62NQWDCfOvzF0Maa11k22yP0Zfc0GZSRYy7s9oslhUlJQ1MNiKGkziwukMG59
k9n7nGmmCuz3kLTcCxHB7mIaxLFwvSDDI2g6qqF7wtiJZ5uXkDZ6UwFFQa7StUrjFrpp8bvx/Oav
d8Gd/9RA/RwK0AUvxuy5T17AwMfo5fmhfTo/QuofdXZ3OzT8XGYN3tNInzqWHWxiZSf/uLemJDkp
GwDIo3UyPQBNoNRm/2tXX2JK1mDeG99e/7D184VZfCmD961qPlY6/dOKtdsMGMfWpa2LlPdlH9ql
RyuuErpOmHgkg5t6Dr5nE+uVI86TuHOwl/5WhakiUzp30XIhv3a6hAoRZ0evNvlJ1jECCui/odII
9rbwanVRrje5vfVs7men4Lt5HAv85wWBUsK1c1x+CLi3c8Ta8Wo2Na11GFV3uN+uBSzIWeb/Z9Zu
9BWuxayF4/k6/imC5ksS0eRo4Wf1c2bsuK0JmN068jeeI4a+HZL6WFYzs3SU6lNq3d0Bq5LBwbYl
ppwqzX0R37MIOk8FeDF5R8b3ROOcsAhyYo6ddlQKYfZ7/ccRf2+LKXvXMrcpgoFLL0m3+8JKw8OR
STH+ZKl9yJWAnMxEkbj/zjoVsM+PzvZ2jbzJVZNzv4dObwzWzPLp6PWRwpnoaW68N0dP/YPxIifM
PjNR7fgJABEtx7SS7hSwZZT7cOu+lMomLuOSQz7z5hwh/JhaBZWZr6XMaxPsmMcMK/P8wE2vFHbE
CG/GeJVwSymsboKNBCzV3LmcCl8MEceM7AdXqaxmJGIEGonrGGaSfJizeYtJijkM+pDqXyeqhkW4
PQznxADW0AG7sSRPS5yt+DwR29Zw9tsZcg3i404sFcGMyOiUIWZi6Gdmt3/eH3XwIONjLQibQNiw
Du2D19i3Nyyn/oGjIzG4mQhYinE6sxNpS1XeNenuW5TSDxvNRrY5NUdilcpQlOQpi/pnFE7L7Qot
tUN9XB9kY/JGjMGYk7C5+Z0gUtdtizKHsQrbMVMReJT1ALGSS+q545TnF+RIBbDurUj90Pe9b9DR
4R72wryVc0IhDkkMuNQ97F2d5p2cZbSza8p6AxjJM/1LEWBciNI+RnbOV9i2v+xTBUolbAyfrNI2
Kf/Vq3J7mIIIMWRUoLkG6ps11tYz7rwJc/ujZdXVc0FLJ5B7vz2gqlHImKUdYSvurvRV3TkRqdw5
yjs6OLOZZpwxgpV/jji8HHgimhNZIN6cQ5Ti5lXJQgzYMOGrRzcprc22jPiwRV2Zpk6tuePyqcYV
cBcFcy7uFeDECSMtyE975F84/h0Mmj7+1IMe92eZzeUorIw9Esm7h84botF25Ra0qbSOc3ld215I
nzRnJP1A1XlZiGpo+DtECFhwmyoSvJrciCb8dNlpgaQALbmfI937izvh3nEQbQZ872QbIP9rbpm1
NGFRwZ0scSbOw0B2SIi587izvJ5t8HTVvCOoecH6RtFguhrRG+9rr6p+lHWrR17R305/T0V8MXqH
2nnZ/8n+6Ct722jc0WSeXjD43A5xN7Xx0r/zqMYcZc6u5g1p60aHNMT2UZ6DXVhBxqKSWrouK6P8
o/+NVJGB6F5kAybdYakuuXbAlQXizDgogZ53qxJvDsYLPJBlJiG5kM57uIuELsF4cvMg5CgXUrlo
iUoX9WYkAf9X+X+ED4oOiNhEVDRpb1x1/bx7+rgFrXZ6deVHVCgiPES0vy0/oBupAXnGh1zi7qJi
eIL0fhq99I5MoBrLsybbTIhVITkdP8LbEtwD7EsmGb+t5v0clxSMyjj18Q6TXORTuUvY5leEUMBZ
mNqmyZOULUwaqF2vxvW4OuafKTeTiwi+yXw3mgZPLE3XZkDAmd0tKMC/jx14rLSRyhtWXApHhFPJ
5SwR9ZetgjV1wjXWV5Yu/4waXo+8nncEsb+0sMiQZ7jiBzYOkZcLhZKCX5VbXWRAbWvcbRAkSTxo
amazRBCZ3VCOY6vVPGPh1ftptO6ZTvV4KPkVE15F9B+dCfgAEZKkh6AbrqYgoxttOTP0uT/gkLJp
Zxq3GtZ5gR9WwARuGjJ8z4P73wWVM0wCGSWM4lk2qxUTr28Pmg1/4uCjBi1ETUPmTrZf2Rf6FA8J
Uz7Nn9E7dPoFyFJ1Lx+TrqAtSIO6D5IxCcXDla1lCyylI+iZ6i3ucxzqpGVuGfCzheFXxK4RD4Ha
iVuuyz/htQCNrIIURoDcy34LqKZekfdaUxcCqXoC3a9RZRrXmcMnGMfYYiYvHf+hTSlzYFU2jHyh
U9uGy9K86hzenelU85LfvZm+F+Ogf/DUV4w9Vc6tMsMXzL6JovnqEkpeZ2vR/E/cu3tim86pNKtF
Gd2iLIlUtnIB9qmH+Eq5PkAw3tP7TqgHO1aPi5ZKdrPrl//qt0ty58V07t72UVKy+vkOIr6Dafsw
dRuKWfYgPeENmLu8M9lrLWzTiK/wAYNeJMD5RLrgddHtE1fwVQasjKRQtWmVjf7w/KUylSAuGhR0
v6EL/XDSTorbWHELc4PaEpHFwETi4v99TVzKhAOV1Tr1oM+Pgk46I4NBvrQZdDUgYn0bG4VLHHcf
SQmAt43Igx2JkJTwUGWh9Drt1o8yZEI2dibAww8xPa7sxgssb6+94oRoSmNOiqDtZqZcQF+Hi1Uq
+z3hbA1++NmPLbR5BnX1E/sojMEHiDx/cpRMglcwW3SA/hRG0+cx2dGffai2W8yu03HiOWqTwE/7
Nwro4jlzODtzXbP0LhEW5iQls/DiUvIHYcRPSHRPnQ+v5v6zzfBpJieAibh9LYBmDMYRdj+1kyKd
uGJt+QGOzrNct1Tw+zkH7T2NaoVqrcdEVWd9bfvjxGGBx+pLBDAlZsf3oPUTOBW78XVwX6hDA6nR
RChG7ED0LgMfEFH1J+H5xSjFHFW6oDFt/l2KqXF8GhHNws3gVol9sA2ncGpipOfRLvQw6pMRRLm4
7Gv4QJWfVAU3/maBVpn8PSkaQmSWemmZz7mqz5CEDe8ICxflGGDLdt5S5OY6735nDeCuRKd2YKGU
Jw8lc2U07wQnOOnX7cc6iIuL/hRxGqPTUP9O7S+c7x0RJ5P2oBrHVQh1AuA1jzXJ3g18Dr8MwSmw
rdOVIfN6VB4S/34T4XlMvzHQALoAf1Q49ZS1OQ/7VGcou1/sgURXbT7WnGw/ImPaJ/ZqemXkVtis
X1Hd3wZyL8Sl9pSvS2/x4XgObzKQpUxlIsyu46KpjuyKI+V63NOPeCKi8D2M+KCBJfMseIbwNnk8
s+EEzymHUklpsnu1Ns6Y5CYgcl8e4SeDskMrkyb2d8lxUBmLMxB5H2N+Mrc4TpKX3HfsH5XXi3cK
XPygRwiBrDxZtP3gJuBYk8lQr5+3J+HYPwGjZP+/RDReb6RO5xER1LCIAK8/yBuvo6613diFMG4B
JYt/ZBL0pzPHw9mT0dEYdJVL79/ylKuTiL+7TQkLEc33XEv9S+or6fDqa11332rPmQStsh2pyvg6
mwz9GN6gwENYMuLtAvl1WY5mavj2tx8zoCOdVyoXtZDvZPZorN1zK8QhSKXRrDXehQkgPBYfm4r+
Oi3vpAIvaZZcgxpGobO71Lwcgyb1dTn0K0RRm1XkXeOMJgFit9SZDq0vkAGqfobCZjlmQywQpxRw
emCvbIeVCxzkSmz74NG4o5ENOFep9W5mD56HPjM3hcraZ/R7APxEIyjkDiLbz9r2uDjKMPonGPHI
m7P7HzeVHAP4QMVoT9dj6sQk7WLLbwIyC1u7vb1Pa5UK5m2X3Sa1P+hxKe6SfylgOXqUPoNSL4SV
Zejq6T2lM6ojirCyFXxO3cZz2IoiNCtAZ6N0Ty0cel8HhppANT9UtwovMMqOFnBvDY60zUnJIETg
WWiGwpvfnvxvUg/65sk4w9enPjusMYlbG4lxys7G1fqvz5TUa8Lg6jrhjlkB90U/BWzRl/MeTCME
hRVHtpb/bSdx2zs6SZRtbPru6AVX+w/42fXTD/W411+ZWapX+RMx2vjWlt7n/SATiqdaZnTJ2jrj
OQlt84GdwaHeHMPbGON1fc1N6ojPOr1kPd2xJu716F5rhzcbI4r01+OfTTyKOYp5u5lUMPHddrjX
XiTRuflxNj2lv1gcQgYvikUUtxOTVYVMmOiM3788bnh/U40oR7SV6NmXXpe3VNdhyd9VttB0vYNZ
3OjFan9KkAze7IlCku8PcBQ0SWf0cQljx3gcNXD1b0GDAoyTnJriBWxZ507N7OwPc0S57ucM5xdu
iprOyPZjfd5yxZGCVCZPR1MgwiQeA5ds6Z/4UPXIOqk6z1IC9Aas0k3MpxVJbPBkVPTHFW518Ovv
quNvxIoAIMOSM8utRNi96mcTYGlvAQGLi7OSOltRk2GiIH++76xRa6ETAFDIXPNqr6YQ9Q9E1/B9
bzi/6K0qSs4Q7YBlrVKaakyIQpBxc4VQxO/gLNHF7++Jxvt/2qESlRJdmj+X1WO7Ii8lyFlfmK1L
yWFA3Ns/dfKHBuYopwSDlKdAYkCRCLlqCHshjuK/l/I+zxuh3xLKcIiraJJU92VV4DFWLKgJoBwL
V6nNM1YhMdNOVme/92HPF91ZK2H5eJmERQ8FJDVD5646VkVTsGDCYYmyQT4Iwc1f9nz+3ceC1dHF
x+ucx5S3k2sAXZUlow9OQlfudP/t4JFA//0PQ5cDq64KEWk6md72e7PzBNTA28khF0c8ecfrFu0R
oJvPieFkbuytfM1xtalX5t6889cEJvBJpaKRwRNnSXnW0xG1aLNUtTXNW6BCBcAdMyp315uIaKaR
6IE9aK0OsNwcc7w3hZfVv/McVoY92eMgkafIecr5DwytQuTqxPYsZkiHW9vVzEdXV7gujZ5nRGHp
K3rD+m6JDmBJuXojRLLmIBc4z7egg/HiY+az/BJ0KvpRVEx2JVkDLU+hP0NGoo0HCQRTvllHvHS7
nb/6O9007VqC1HFxJgVlocxAxjPdVoeEBQzLVXHauSPSksj5TPO9Bd3QqJ+HS9KbdgVrOWFdVqwP
ddjEWiy/GUv5dPsxn8TW9SWsruKOvDViHd5NtiDvLFqxPZD+mK5FQujUtpDmcsOA0HSQzl/DIcWu
zMnYTekir3g9STOccgevUX/vpRCbbPYKdr/LmzZ4OEvqgzA/hPjdpqx2UXhB+Dqs7NLsaLl4P5+/
PLJWg9Jzh7miXC7OtBaLqbdopyKQHCQVlQlj7bC2GaykYcG2YxJe1HG6Lejpa6Z0NY2IzTfh2vN+
qCzbYRNwjl0MxBQdMS89WFSVVJDoIARkkO0iO+VN/ebtpw10UWT95FAjkJQ+krYqRtzTuiesNDWb
mRC4De6o6n0t7WieizdX7cKBSbN5DzKBUC5yta6tMRorTxyoBMPAWL1soIuVYphtm5LT1QIStAQV
F6RYfQePReUj+vOXuXBmBIWhTexTvS9UbrQ96c6+Qli8ENob6QqfQIQ2cVnmV+6pCKPupf/U2N8p
6AVqmRPwEtyW2ZHiaS9cY1yUWfp3lGrmkxi2qJXXN2oTotXgUR4s2GUuNKw1xz6iAcmbQ5lyDPeZ
sCqSZAYiaA1OjKuL+h+urgQMF4sWs6fP0D1c7eh89Bbh01v5JIWiUf249sHL1DSMVgHuT4qGzv2w
0sC9Owg0L/HOY6lHQmc0GHKzLbXI8HK9gHqly+neYePRGX4dXiYuDQUAkkizyzWCVk7Lt65npibZ
BLxzBfPDFy2n+ThinRoOAl03A87Q7MD8szKUl8oBoUWnbid4DNPlh5ICtG4A5dNgKpFCVRqrPTXc
vK4v+kOEMiQTEJfGoy/U1KebnWk9P+wkccFyTkBRbdtV1cS1o9K19O5AIiWhwbusYN6K0zLIfqrk
THv0mzirLKERunj3v655b3FGBWfSlXbKHKnZSkzJ53+dqOHlkMk7sYQPOOpe2f8knyJBQdvlyYAl
mk6TaAGMRJXQ4LgiwCgv1xEfIkJiE8VHtiv+SzDoBNT9pzEpnJh6OZZrIymbFdNxSt+mnTiPdJyT
iQ0mJ7UxNFNAnSpr1v446EUkEtVkkpUhXMiGRzH2pDdqT6s1NOSJxyuFt6KglYXmrUoFP8Rq7/6I
Zsgcp42j/SpXVFn7cROlppeeyJ3uPiFa3dPFAVRS1lt5pz47xfPtPKaPhoq56eDrUsAZwJ3Jjxih
Z1sxx8q9FDplyteK7syLzb0Bqifl5sgrtvPr9iaeAsS8MBW9FB2SBc6kpiPCOqIQ8OA7+3GbtDZn
i4sN8VqNq0hDb6QPNJbWPT2vCmDyNV2wOZXoC1pehz+QZ33wIEfMeIg8TsZtNa3jhWwPab7+lWsO
Q0eBKmjFDV8/WE2E23sIKgSF6vRwtGw4U/Yefh1zHBhCOT4kMgMLPFQMxnkk4DiQ3S6ck2AXwuPl
9m2v5vT8NtnFZFsxX+GEA01vTbAXVXSsSVQKKTeYSxtAuofFKrdk6pNRjqkFoAAbUPHY3Yg+Sc/S
6e+yb5Y5JABBXKlU6N6sAsx4VjvwjhHQu0WFt/lLWJCDHyjx9eWAmKHI+kQOQlFv078P0BGlBeaA
aSjxzj7jddw0cXZ5pSVfhcDwnpUoqyDlGXuyTWEktZjIvKC1wNseXH6ubArBrsr4bJeovmpO0rGa
fbnXAvRJNVkYPu9sCZlGeiNFJEX6whafd/+SmGM3oM4EozG3Fw6UqNxV7kOiQzHMGkxQA7EAgT23
us8CkT+l5fCli2htwt1/ftI4z7IyCIy0eqyX30A2TYNIi4sqRzWEekeuae63p5Uxg9VxZW/Unoz6
EAJvY/A0LxVaUS4GRgcG1EySipO7MGn6HsB02pMcA+FR9IbeBR9EmSEY6g0h+/JgjKYoCcQ+pvEy
SPollycY6QrCy8O+XltDOQtAg2G5EUUpzTJvAqBP04roPwbSn3gwaqFcgnZCY76GGxOZZsRyvBpo
uwmAEXwqsxBc+mQ9cR2TXc3zyln+wfCQsZkQxZJIJYCOMnDXlNwOImz8CI/995cTEx8mMjOqGcwd
GQ7CFNg+fU9wTh9MFxlXTxeQVCiPAD5aeLZY2YTsQ3S/P2uF4Zb6wGnip25WzVqKNQze+zNdHh5v
ClGhKHm5zp9Wl3891DjUctsYNlFwYFyMpBgjSiZf8c/kNbof5AhZ63dgERb/8D842e6zi8ymGLT2
APYrbhuvh4qjjrKxSsEW1VGKJo9A2v+RvLgqQ5K6G82k0wlhyXIwO5R4tLYdFsdMOhrXpBH1hBbM
Edi9miHunCX5GL2pl+A0RhAp6CY2snHAFC0uhBkDz9ekJPsloyUzmIqNRwuJmOSLGlOTb3HPqtr7
lZNtq5+63r7hhwMuEE8u0CdxhVBep/tU6CdQxUKn+lGUIlWTBRILMvjfGIHfYzoUFF1Bhz6e/TBF
WLpazDZVkyZJj17UaUpWhutkJ+Qv2FU2wMU7boF4uCzcLeEve2pB/xYEg2vF8uW2i+4Fd1yXZ1Jx
8IYJWhx4EmiMtn/76leaQLjzq2Xaga/N1qsmewRbyYR23WgXIiKQ3L1t0NiaVQBR6uWAruuM6jA/
oP3X0nbGpHePDKnytxo3EOqxpZNVYfnPSbTzMN28fdUM6zyZC/2abVR4l0Ay3EtCn5GHFhZir4T1
Izi6Tmg6+NZZMLCkQ//OJIK6IaP0MW0JL42+jH6a8UZnt6a6PN88U5heauk9hpxLblcpUqnatQtI
zmKHUbgqByF5M1XfCJvQl8H+BsnvJ3/SSH6yLreV/20+QSNpgEeTybbLPXDalLnZEgAjw5YfsXVW
X4TPx3+Q0y+y92j8xRqxwjNSOgVoB0CF0XW/U7ZEd9UfapHACwORu09GluIbrJjCj2crcmEWnQ4z
T4md+y+Lq4mRaa0yP+N53Ow3gSbqXlzJ00s08agt/nfwtKDtPE9+uogYeq9AjJ/Nl5DoKspsdj+T
TsPHtABiXJLsaBKn3LQykNDEmWDBu4xTjNI9ta5ZlX8PG5iJnD7xZ2bx94LAW+4wHLMhscfr9hDj
vPw7ylZrm5gZgJHbrbPRE56X5dVG1k1Bh7DBGTXOAhFB1GmtSrLi1CaFme7CVQ0XoM2gyt5Id4Nb
rjbwYOBeaI+JUU2Lur7dEEfUOxcqi0dyBSnXxw7OX3EUx0ni+ow69DfTQSG5vPUzxm1EywQ0LeVv
8tCcP5omxTm7t16xIDTji2abTRPOX9I4xL2HDXQoLTpduqvOTMscF/67DSe8EMxjI7Dq4YKKGFxr
N4D9AFJQgiLd+W/e/nH53zjlIs8EHPDSvmhZBkaYQgv3mf+rQVubzGhEnkqWqk8Tp/vvAkZXi5XC
gaQN4Hw9T7H19VZwbXG9FO7wRtO4477A6TFAz0e6WnABpzSRUTU3MSGefdNuZwvA/kKFfnN0GNsZ
3zxe1QEuEiWloNcl4zINEfKj9SFpHA1rPD0msGZCcHj0BMArLC88tAjdd2NiGAUnDZKKqGihqy4T
fFKsdU9C/EgokBc/+yK7S9Do4rswMpBjfW5wL9VpbAuNy0EpIuxUH/tNAqQY3rqllmnxeaT/Znd1
KI02DDcub0/uZpkenGr5M1Z26UC7ADc5/Q6OupKkM65YuekWq634DViRsVLgfJSdneYsL+cS7n3B
XpttLqO6lYlljBVxwg2byNrsahCvQCeXLqmE12jw4B8AeYGilS8mo2lsdyIi19fBz0ExP19wOUtl
yokZqN5oJWgmrT8KGek3BK5XM/Q9y7r0HqRrYnFzYHyT6uK3yJL3uOXhINICYPg4ytXcyqSJwt7r
ebR/1eTCR8NMUjAcSwdLHrWGxd/cfdn4aeDkMg6pC6dmh32kdxds3dgFUPKnLu5brNBVbrjSkYvj
BGojbOgxkkD5hnAaLuYS917qhgu4hXJLVaoGLfUP4QMh+KmHo/QFn8Dqa/f8pWiBMihLgnakO9lq
jhE9jP8bNxopN9Hsg43XMtUcZgxAbmgbGrgXOVClxSP3kNnTdgpdfRK/4vWoCF0vGAOprT7+QIvQ
rN2ljimJV0qOt5No7q/GypFP4iRJEUGLxg+Eqpu+1gMxxf9p4n/tYBhSGBDH6UTBdYAQh80L296J
b/AxHcm8TgdlJikgf5TieTI3m2fGe9pPjAJaZTn4o6zeOEO/jXweZ4Hvbf5jtlaTJZftGxNdnK7r
XCbTsxiSVdx9CRuAoOtU/LQM6KxTlpczdkJVYjBhKzqhHM2ZXvxLl60DDqeiYlKQQVfQBpbQ6n3b
JYWrdDG+fJIm+xZaSdZK59LznsGMCpXf4O6vUPL9L9hSicW3UP8+OvK1ysUEtrXd4SvlWjj0NVfR
++nw1YFF9PeWjwvrq+PSWzXK1vCNT5UCMqsTVOv2/Snfor+ZHMcEGGbVUBsx9DGm8m3jSEVKoOHF
cjNATtahpQyJEt03IfBU0xpEJK+m92TJNWBtLRBS72EZ+BbnzHMb+ptETe4PoxxU39m8QdohdU2O
YSRP7lCyWcfE8JyjvChy1FDXJpmGqYl2a0kEVP8hnUNgKEJDWm0DVXNPQQwQeSuQlMPK5gFnzLtj
GgEl8gyIWMY0KS7qs/oo0dSp7YnWyo8Fkh/LFKBcY164JI0iD8TkCaxm41LzS0qYAdpLMj6msxF1
ujgwIwg2yyqffz2efCxTwU3N6q+BnSEOBRYwPEV4WP0hio7sq7WidvKU8hp++LEiVCGzH6f0ZgvZ
qP2tAgsJmH8Jy8XGQcxNrGeiT/xC0aKPNrb0SgwWRawr7MS3Y05HoD4pHbKL7OR7BBATvOjdwsP2
nZp0hU+VJgX4vXA19vUN3TFhN/MkZYDUNbHVPGgShLtynreW5yDg8p2YkaDJOT//STZ0xCWfBYxO
Tjj+AesfcHy7y6j6Cbv06KTzjMFI73lXUFnYtE+IFtxiDrh43a9cWSiQOGSkwuxsru/2F8k8JICs
dMVWDWAVsFO6sWpVNfyE2Q44VwSkaaeYSoKtKwxMikpcNN4VIEpBb8hd14kp24dnI0qxUyVTxrzS
g/W1AApzf41sHhAUFZbGYCDv+YNIrFZ9ishvGPso6Wdb3IPyqXoWMAAQ2N1D9SwEYlErUrepFTfF
Hjs3OE8XuGilD0M8bclTatFBrKznEAQnrADJyHvoutRrN6lnuN77fYCbCCL9jaFmWvXwVP2DgGsz
Y2Vhw937F1TB0kgtCBlTmSMqvhsEi83FbFjtZXNtpVT1xG4HqlccUBsjhT3RJk+B00o1L1mME2AJ
YeF2Djxdofszb3/UHPzSgmK35QBr3NMYACeijFDBHqdLIiJl6mQAo4aYVnHuEkSkIaPIYICWEM5N
E3q6tP0Xlz8tOlRqMXRgOdI4Cx2LZxbNj4VXqnjWcrcYlEt4fzc6GhRw9RN1N+gQDjvbhFj9TbM6
6gxanQu30LVB6nu4DunNN7XIOw6ihrQ8w/wgIdqk3vCL0c9FEgGo7eQXVeKR6B9kNMLiSaDe+qUz
HOXJBEvTjDLMtnl6PBObOIVvjjXjpsiTJkDTloHv2s2JicaJprrWvIWS97idYo4qNBey94DOIBaX
E2d9E14w63OH5E8+12/kEeiCcoCSlHKCBs1dCZvVMnoSWU3cHb6nahMQSrrlzqVWWIKeSWDi3hiW
aaQVgVegWvVAKTF89KBZYcR34Is/rteuGHKLI3x5FuvI4AfIUvmJkf6VtGFng6rYijy4Tzq3Me8X
scdbK/2tTyPyWKIdnbgauaEpeTGVED7xbtwxglQnmXDTVzjbgpSm2k6XSbdNnmqUPZkU3ZSobq32
FDjZ/7b6j5TKyva2e8uS+JA1HaBzfoFwsW+Bhu/wy8smFMsrfqnRYmgjxiet5XBR5EYsNf3YoRLI
J4AhNV/Sp7VpeVIHfmICSL4/sMQZRX+TWVHPIzNAgzdvqOiCpEvVlR7XIFp602r5mPdheX0kph5Z
1upYQ+EKucDIa1qpIjPFfczbLmbLeQcPAbnWR7SxBdg6UMFwvV2AKr/2mIeZWEGfVL93zGxkDJgD
hk6kX+4ZDK+Xj7UovIxzaRqqy3Jtde/MM+Iy3YmQhuspYnCrKzcHCSDVSkbj61eaO7LyfMwvGpcD
gdpLiw1OsAmnCrJbiS1qJGXuCor++3Wqhjc6AWxqtHL8lx+BFVq8UUT35+WSnhVNCWfvZEPbKY5p
Y1/q9d04SayFjHhn7cbZU8ftKPIwWo35e3TNGjv+BL1J2og7LFKj7RlGsghSWvwZJE59oCbIs1wi
2JBccybiVPdLO0lXMob0yzRDvncUV6RRTDmhQ5KFLL6b3H9fl05jcWSejnDyhYuNS7EljGt9Ziqm
l4XgLKkVbLpuEchF1ROgCLfkgHotxqiVqflW6x/zvrLO8BqCUIj+fWse9gjUL7VlfYqCQh/R8Udn
AD/GL4wRah7f7EndfGob4lfI32PbPb8VjJWF5f4zKABGvigNdvAyB66CODsymdSDvnn/oh9HeDca
q0LWRBu3pSB/Ez8jn2UAv5SiD2z9S2YdDIE+4XQD0H3mI46Z6aM5PdYG49dLNdaK3vt3gUcw04lS
GImC7/K01bXucrIISudxf32YxOgd+zPRJkSkSFb7A1RiPdLV37m6cKMqDbCtMX3MqgTu7r8j6sI2
facOkPI9cGOJbP49P2N+Y8WfvC97t3v21zkPiDuMJavHt3YX42npLW6+KDulEEvi08Ei4J8Zxzd4
bnQk2JHBfnVI1SAI/e6srM083bqduujm/oWZ8WBej+Zob+nwQGOV5DXT2sFICXsb+EbQvnfWvC+c
E+N4U/7859nsvroNmHxk+x7fI26Ndsi2Qa5/s4EV0EArbvO5QYgiUe9zq+uSP7ap752R2QH0IWiu
yAUmzABh1nqpPZ8yogmHvY1PJHd9LIFBI5reSd6StGOwPZx79Wi6b+ZGNjx4Vmx+9z3DedA6TCf/
UNQ2FSb77vpfAQUtOHgSj82quS5S8e0Kf2GwuTfDtXIz6ViOl37pOiAzOH5Q5Wbfh078wfiLHIWI
cy2RxEFH4KEkDn4XvZ3iRChzgYqk7F0LJFPLo9Et/ME011YjzfXvd8kJEW6saH9lKH7Nj+7aBi45
dnMasX/g+abuSbG1fRHIbJDFSxkWJPC9xaM1V/LJQ686HW0tgsiG48QARipdyvZGMoONWNvaky5I
TOeP2+yyRxXuoOpKiiVDNmTtdsAhEwmqMhLwX+zPimkh+wjWw8mOeIHfwW+ugQH7P3NkP3yEXl3k
DjBA5Pdb0fUklpi/HYP9ZDI0S9un8OyFo8+4RYWJGL35QcQwPeBGgbeLjrpfs7C/ijtiY+7l7O0+
/z8RY3SyXScHGaBkYiP+NZmxaznVgRG0uA5uuQFFjmijPBAZ6HjnC6y80qeCB5G6P7K11jnlSoNe
m6lvQ/889ml0YCefE8JjbLWVGs5z29BVsVhq/GLhMIOMIWNKNQr92w5OXhsp4ITOk92sga/5c0Ay
06D61B7NkKeXOsJjUP4TZbngFqy6QWHWU/QIYfKVF6mhjPdphcofo02qLHvntoV9b1J0dzpXpVkw
C1Q1IaH4vhWeHSPqxa/LZ1kEzz5p7ULYtiLCpkNDti+b6YNUJoZlaGY6/GDwZ412xWLmL/XEPHDa
WsvcDOibIaAx947ylPNOGpGUXxPue+rU439vU5uA2k92J0q7z+qrCnspKrGMQELunvESYtErfv6Z
wZSDwqzErTfrRQjCPdJVmZu5QzSFwUPcJJ9Q2Mhzmy8ezk51/9ysp9wNOaEfEekips77pgJxtQDJ
qqydczMuU+5/CJwpRdtWIpXS+tFT04d8CwmP0jzSg2KnTe6VUnl240lATd4JtiVr5whkpWdQVaNI
xmBzLQ/W/RivHXlKUHFxfze/FN+scq/eRkXnZpf1vU1H6yHhAO0kbr9bTMIXN7Afxj5WrR6/hgLh
bJhL8Uj0RPA5gkUaITL5fsKZBrFCg1MfMCs8e4x31Ds1mKwpytBxEwNx9MusF8rG11jzwl8a8Ww6
T3qc9lBVdkV5i32ZW4ZjbzGdAq1J1udMajbII7UiQf8O5OxKdETkdOgWgOTKp4rcwZCko1c5V2AT
YbBLWjMn2MCVoxxmEGpJX6AFvV//v0O+8ajeBa45qaxST+GZ4m/scU49QaOiNR+geCQiXbaPk1mE
oTlugZe/LXCPGOWqH9lIin6hd24EX6xl7MslgSxo+jhF7RwXfqF0ltbR02pKiDGyWrIoCuA2dmz2
bLQYejnVax3YRwRVLdTRMOfMWXEbQjKePab5EISGLMpXDjsUdHm8nSN18Nb0GYPEeUV0NUC5Y5qM
JuTHG7yA8tXJAer/DWb2b6qRMNisSS2ja0oS4BeuEk+P4ENiS25CbwtNpJPUcczZvu3uSLqzUOcU
86/cFTbCBQvUY+1MYQCIp/3xy7SbPmzh1rkXr1t+raHfV6bPec/Va3e+FaUKouXj0aAgnoN7OpR0
FEFeZyVMZ/aeoD/s/Va+6Qg/CIaw2XFWdFBN9xtNMBn+XIRvg/1eEp6J+nxl21NFihX/SYQVyrTD
AVx+hG9ZiWR2xVJVOi0EejiOGcpQnQnJvR7ZiOuIUvkab6Hffz1e3Zou1ZDNb2Y+PiQOYBjI7OeV
imQARlQ4HV1ETVdWqyF6Ud6OBloNlNoxfH4P9ihV8GSwg/E07l6k4gjHs6r0lBPcmfn2pRnrQQrK
PwVVBp4UEmiROw5DBRwJEm/lmOBTjawxZ8P9/KNJYgnnMpl+1Qb4MhCyfesaKR40E4M27Uf/h1cO
7CpHnBSh/b6JqUFofp1GGQ4THdxpk6fhWX1Ilhtxk6Y+zl9TPn9w0VxNJdXGKiFUkJZmXmcTXe1V
KLSsQV4fH8Ls7do8yoeoYCUfXfbIvQ4bl43ZQHslnCI65jqCoirbzzjluISDXY2vtLI0VxuF+avq
Gp780KJNyrImpEyoSVRoabKE5g2sJ5trpjUxZr8R7EWSEVtTu8CwP5PAqDL7oSwN4oWKgY5B5Jaj
4U4sEsR3eMHi6R+7s+0SOtmRPnarr7+7oL4Vt2wTu9uBbpVeInwPJpdJWmE4+YT6zWU0f75Drl3a
nvseiJk0LJjHvLscyO4ywlV8BMMh2VwdvPRiJWzSBTL58sTJKCNn+n9nxp3pM3DGPBP8trYi0VWx
oJsuev8j1uTZ7HOmOowTHlcFRj+AKTPJR1rPNQ6xuFpA04dOPaZMm0c5HhAiEs1gaDlOK8bVXEpn
t3MjkGeOImlANMOkcSTxp3V7kkwkEwBL8M2RMevtByuhI6pvqwMz2Dk3R7KSKao4lpNMltGB23le
wwCKm/uXPGK+rVIeQb+lk5C/s9wq+umVmN2wqIQIwCGUnj2vsr0nOk8WbGwcitkXUuIdI0qbL0U5
1laOjzluPpPui6nDUPsqkFE9iUhX80uo98f5zLFaoaCar74hnj+adICudEWMU7VyJqzf8kwReeIt
VzbWrtNk2MSzjfV0B1THWFgUG6Gz5Clbhvv4dLNms0ukrgeTvJqvvDwF3E1qvs8jUM41g3D9OR9c
/hfVtoS067c6P0QUEXVKEJEPMi6tL5GKt/crOjivJOKj3GySSggF2KuIn4+jrUwzFl439MvLy9XK
q25THBNCbJHhqA2rGVOzaswonS5KwO5x/rHd4x3NWkZkRPmXHQ6alhjW2D+Jk08GBf8uIlHOQKdI
a6I8VBCtyags6Ydu7nhaCPZUJrmMf5DetU7uPSdKXgz+a214EmQzKxFw68X+JfxmZhwCXzYez5L3
Jhh/1PRk3DnN1ofWwibjn4KcuzQ1KY7lYVTdrJDP30kvM4JjEiTauozWHnJkcWqboVStnMWEAOqv
NV4zn2QY75PQvvq9VUOzGFjir7B2kMqvzTo4tCrjTUum0kCZqu2YSX4RbbUqmGNf6R5y2ByHwlT6
oi2eDKdzCtJZd8XCtTCZHKsoGOwlDoZmCmzjdNgSpYXJ9psjC51eZOapRjrUgIQvF6FnlgW8TH+Z
dEtoYOSifxO/kAwuVNn+1hJS04X6JVAAlqEfkc8YNceoBsCnJIni+39hFyNjfmqSomFbWDA6aTJk
sx6g2trQWziPvAtem+kfcR+xdBorf2tFKa7zQZtMPp1wdWrncsPBriKAOf+/34Qw1oRFXcL5ah8V
CjToV9JMfLKvFucElxSEl86r6wOUfgmnmYext9watWcvRAdp63FYdaSbqAF3pr1lg3zKzw6Ujp1a
gyoregUlIfQVvoacYGe5Gpt5aYgAi4EXwAukYqX9FE3utuwq8rhgS/XqVJbLq/oB8qWOUXm2/hCc
VywgrRUUPsODqcQn2vkqUAOps7MzEK7WoQcWBTdyeFT+EjdHX/ngHOjn1hbvJL+HBvZJ0cSCb1tf
H+MsRcJ2H0nqcrN46s2qH65ecqH4DDJfT+3vUpx/A1ieRHfQYOwt5ISTaQX3iWgaMD9oDzicT2pd
ZTLqmyAw49GnOQ7wECAWEBLOYnMamtRlkhKNy90/fNKV9DMFbbiqHbTIoSENm8FByO8apB4adc8j
dhpwrYZFoMYN+CSimHM5RJdfl0I8x7uH2TRB4nLOIrx2KHJPUgQtspxpTmDGGRxqbNBgUJ46zoEt
Z/GAEHH9Ip099HT1oYdMB2UlqjyOxSgW/V41SaIsQi0uePvcIQZSUp6zFE3SRK+FNjl1yDRCGyU/
z/wCs93LhnLnDSOEFOdspz22n61+4vtg5E3hpO0LuOwNo8liPQWV71edj15sE7i6IFZb2wNV7Us9
lKBBfG+9q9eKD0BQNiCuMzSnsxdJZSCffkC5OVqcTDomU+A9927z5Sip3pz7xp/ot8tOpchTRnJ+
yu1OWQEA11g3IHqLOb42wQ6AIKs9s1t/D4I8EnwJ0s4/Z2uW1gBwSaUgqXKWoU4FuCMx4XzC58tn
wmZvIEUrmal5bmDUBOc4N44oCv4ZKS23W1qON11g/ZiOGlCIxBf/AiaVkVuFkyH9zm2bBJmWBo4p
U59eDjdcPgu+f6whbW0AUcXOt7RzL/XunvMVeAoXdFFhFuaRb3mjo4g5e9YeTiTaJYx8l/NryK/h
N8/l01yawKBh5Hb84+DUwFmOEO2rE1nRUqzSgPkUn4BdKVDmByqSs9wUrXAp2+9OiLWDJ6d62dqU
sVVHlMhRla1BzbWPh5Zytieql6pzvrd2hrxlzsheCBit1hSvBXBIkkAoY9sIg0EzyCWy9fZ6namF
XRS0gQTrNtsClb14oUWN+WiZzO06O7AO6A9DxWMBmDtKYtVpW+hhaytBnTZh/wxSTd6w1Y1vEog8
5rGfLo7qvelgyPhPnU64tRJxu/YLhrM1OvJrtPPqaNU1QHcG27VdnTTeMENYiXJTwR/1BCkbttto
3iHvYlPNmKSGZKLxWXGaWgd3iAzSozdzMAZUSsZGYDtHrIpPdebQNQ+Y8XftVTPR4J+6qNmYg+Ac
WFFMJk94M3Hv5oH9NNG/a80bez3eEKHFSX6yZXY92oxb2zClgczgmLaMKgvIM6d92JDX5Z47bBgq
sQKXARAIsUzSKHhTF9bKLoAsuO42OY8EyohWPU6d7sssRp0lRqjwOZQMxeo3Jrm0OKLzFOIQD0dP
Eo1DFjajhoLsmil8VnmFGayxavzSQi7Zahm7DuBUl85f0/OzFuJnqHYDzIircOIyJhJTYUSSOd0j
OZKlRNgX4AwZIA3+vzlBabPmtYr63zjIsP27fJddJlcL7UTucpLpR+juovKYm7Z9hieDYZdMbQFp
MrGb2cC6wHQZrsuyrBaV73TuCDrIID/3q8TizegKQhBibolRo6q8VpVjEKpvKBRfgOgLuj9a1Ttn
HIY91cGgocIV1BUEpZxBe55GNnFXrVvWIOIzBlC2zh93a9zvSP2fv2bNOPDcpKpl/WeuUs8GDb1E
GFfXo/R5LDgErDtuHfqzyd/hrqFFILhRBlYLY3RcT2pxaW1i2ojMZziIsvwRDy9Pa8t5hyIKplar
LRQH4YQsA7ZUD7vDYn65NBI53YlZ2KozT6ptV+HO/fmiSYmwxGIjxqipvO6se/dVWL4X4yea8FDx
XIw9ioYwoHradL9MER6ZVKO40ft5M/MUtuLJSmu4lTXzvEFtaFiZn1R/MdUDPn0+Zq4TfgiM4hqf
t0haFRsLNVOWBa/BvIfN6hXY12og9AGYHWOvRmbvg9AIJuh3NDlMOuBQUfaS5xQ5zKJyPGAh+K5C
4xLItzlM71WJzMuHjj0vOd9y12YT/jvxcziMTaTs0yzO5jN4AihhihhX5afMncqifVl+zZ2UCwqB
BFgTFvTsAalWMSe3CDzumTELE25pQAv4o7UndC5VyMadZdWTW4YrAStsGVXgbMzmkL4M5xADkUHq
nmqrhN2muB4jpMACbqm1ZWmRXmhdtI07m0fECjwbgTJvvoXOWKMC5ekMCn2OOn+i09JNbqO9Qhak
LSjSDhVMjTL8huVRoJJ4jHFpJmLglAS/Lb0M4UDUmWoP76c5hoNAbz+hpKWajMHLvW8nDZgOSHkm
ozQ900s2/qwV7Nikr2IMtRAeh+P0RS2vB/g4avmbJrM5oz0k1SgQEU3ehGBhF4NPED0u0lc1gyzT
YKrQyEMFNxK9C6CHuGgpTZuPFsElf+zMOH13DY2fs+b41yxuNHXflh9b8grZYzkNKsyd3h7sLB9S
WVs1NIRL3Hs791U79k3U12ChGjOJsk3FqYAe+YbWJfwxP4HTs4QwsFORwi2dX4MxMdWAllsBWQFt
/iakoCv/KgA5wxYvvzQS1GRZZYau3J1FSEiUu3AzWobEBk8Pat/4tqMELCJg0/PTiUBn/sgIExZV
/TFb12WzT14Nqo0l8QOX05yw/kOSXCliwdtLOsk9OGg+VM6T2wIdO6PWBaz4ZSgCdR8hOPfVMNAx
YYTa5Iin4N7/yYhhlJ7U9N3r9TVyt7bcC2ethXuj3ORpWTZm8brOC0b94ZfUvXmvjX624dXDLv4c
gjIvoSOvqzCzZGNsZBnICnEmo2fYxVmWF6I2X4GakS5/EPLT4FRVf77HPIF8thi50Yr4qinK1qbm
sCo7+GiNpsELeSWUPFIhJAqnmZ4tdPbRQUN7deVpMR8JoJUZW4E/Qyla3w5BVv1T8ya3RMelNUbH
Ze10QUf6C3Esee4ZHg1MtRZogYfTnFYx+IfyOlXfdtfaxfm2Aoh+nF09VE8HG1a40c+eMJ3JrhUR
hO9p94dHxaFeiWOjX0kIunpTZeMdCUTMsaXsmaEFcIEfSQNQDD2fl4bwk29gsYIaxqyW7Y/KqvsM
2MzD0vY7FfG84fIyIvK+vHa12tj92zzCwN+5ieq8yeZHdQp9H3Ls3ybKH0Y/i1QRbQfQIDjNVK4I
h7MucvfWc5CiFjebqxalzP49tdHcYrcKce+srEIioLpJGCn8xKTdJOgaDfqdMR473Q4wHJvcoLHn
ho7IlPMdaQ6UHzczJL6nP2+06yvBSQfbUIqXP9hzCrnZ+2Dj0Fz9MFVuV9ofv+VkZ+fFHWcUhlwP
xys9wMgl6JCBSvdQnuospLZU5+EqqGPAG3MVC/0WZc0t7R0luB4f2I3xLB1f0HiRsDGKsj1ykP8z
oRQfTsmsBnoBY6H3Kc8T7HBMEngTr6MbvQ85+m2ZBux3AizgJaVce76eyDfMQHOXLoqahcA6Q9VN
/9HsH3NYJ/XFCafo1NTf6mgLfNAkEs+5z3ujFqzkkdoXFpbs8We3e5OivtKYXoQ/G+W5QDRfJW3/
jOSZph/0AomZ7UE6wqEtzPsRlmyMafc8ErQA8zb7vms1Kson/4G8oYN1pE/6ggwlG1i4P8fmFKQp
QWO2zJ9vq17ZgWD7dNm4eHKm8R2yu+AeuN+XsO6ZPkypbAk9iq5+tfSYGx37qCMNOgNeeqxnJP8l
THFbk6RseMsIY9S3GHQ6c/HupEExEgh8nrZ5ugSRERp2U6Od8+htcksC7es1xbyltRJb8Ox9/x8s
mT7xFYvZjDfEnoLQiTZEvGUPGZhk0SLsgYh/bHLjw695H59P+JmMcfwlnnzS/GXWABFTCWysJKbB
2gHFY3VRbdG2KX4aPCL4b2qs7VgGdVM8DE9K6iTsjzixFYPaD8AonYsrBkqGVBCVdVbNaDR5xvNq
ruK7piYSPYvHaAHhQYbHUvXqJfrN4MNMQ3D8EWVwFH3oarLxmcjtMqcIMcLIpTt99Ka3ZHL3w4lE
j+LSjhLaehXdoNA7GKWDUp7chxC2skaEzM8kaygfKtaPkZZCEP9wD/9pc5YmYK1eAo40aT71EG4t
/pFm58uufHyN9cn3dLHnTcFgMdRxR1lvCnMQRcs/QPix5L2I/m81DoWj1x8xYH3rdsVStTXdKKYS
439OMYxfqFaJM8ZSXWkhBOrW/ZUk2Hstw1souVbK4fYHL2YlbIKoIXVu574bcVDX/6QADwYJY9V5
YzeKIT8Zx8dUHPA0pigyDWYRJXeqq16scDiUDHj2eQocJ5rtg1fi1Di0AKYX3nHoMIgNDuhO2of+
Vepxc+UnDVPTJQrFQDF8ndNJj41+TvOy11s0kOpQfI7LrTtv+8cbBEe7b83H7q0leUBdATFVLdk3
29ve2qt4dRh+EKTi0rVaDyEZUeyY1Q9YYJm8fWgdUKDy9r7WIjdK3nHTB2ipHtpRfghFBdqbHWuL
7N3WJ0hC02QJdXUAMtDqJBjGx6sewQAFwRuKDa/dLbtWoQ4WEI4IKswoxSCKv8Hg+fkDJIE4N5JX
fdQ6z+xO/Lc8BISvLHxwEQdFtwwN2vCe+WCaUn0JJgLcJvKvr7DPX4K7LeFwb0J9r+Cl3T8m8A/L
ecR2/IpYlY2CfMjUiIpgNDcEgsc9AObynmNtMCm8P5ElGdm8mg7E36fSeH4YJX+foMNL/7jX5je7
cyf3iiI1lyND0QLphdooktgV71XA+DhGGFPWAYxc57qssgqid8uK6Yc9Pj3kONEqL5Ot4KRSojcl
ckS5obSkJGWE1SKNOA+gRpIspLVWoZpIoGHVSvX210EcKBQRoI18U/Lmmp4BPrYzLgsybmciLMgS
xOly66Ej7b7bxYECdN+dyGItQsfCaSIaeUeL3jh7sQ942yv/G/kTpSKnadjDI6+qyJjf+YpiPcTH
w+huEAhthiDu3ruU+uk4ylja7FvAnnaicz4mcQ9seFQKhta8tem/A876sXFf4F/I9/UaMzsd9/4H
tP/zF2gIkPucODw4Sj1GDPaja3ax+bGKDteZLPtpUyszzY96+A7Hw6FSp8f5VAFZKCUCx3eJHj1y
F9pl5dYtxzBsyd5EioAMthAahYOqP0NNmiWGWya2S7TkxyQzTUc0you6GIG5cUyQ579BC4k6afTk
20bSjv8qdjabLbqwls24wANF0GZj4FHiwRv7zCbrtuzQCd36lswZF7k/7mP7pnyrGAKCOmsdr4O0
VMIFSPvQGd7dDvO1bePb5bqFDyZVVXdtzUQHg5VJWT9nQRM2Dnuika5gZts8pnqhF5B5ruey7Vzi
1BWiquGT12xKKH9QigcV8qFsv2C54kyDQBQ9A1FDPd0GpMNCl/naxDL2pPudn7AH+PME8zFREotW
4ZI+HXIkL0wlV99lniR4niyf1dEERRAYOBGIWw8HhdqTWoTvQViO+EPeTqF0w90IglNEJpu8FMyG
jb9kOU3PRbsTb/+DEd7LoC/3AvpsrkYJYfE53/rF0EELemeuqYHGmweXKEuJCZVeUXYcqcqe2/Jc
wq8JL64+k23BiTSpG2LPMKD6Bwhhl02lSxO0hi+UKaaM2SFqC75HpA550lTtW7ZPNERX5u4yzgYz
CWljzIMwbBc70XxDquW/ZvqfjjM7+SC0B7W5C0xwvfzfwSviSYqIMqMx/zQItPHIJHHwJi8GH9F/
l1zWOe2c+s2goBDugGraJwC2eo/FuTFNPLwTtckyc+WfSwM0kfD9pWPhWO4lGy6FwBncnafx3Q4F
0p4buZtHiLZ6FrdT90fKvgHxbsD5D7b2wnv8TdYe5QBQFxa2DoD54TXAzI6NMnBIyGZ9PNhgcVJW
xTQKkMaow7AbHOmdyvxmTXnZP92Oi07NGZCigeKYnbS3zqEzaNqhmDgRSCII6swSEvf7xAT/dHXp
xldZucZGuOymEgKsekL6DrXHicfYuHDKZ902UHXB7B3caJnSbf4D5b9eIsQh+HT3GHWzcSt0cHYQ
rF9JZzPiCNPV/BDkbl80bAqBz/8Dh/qDwKdasT2Pu9MTiQTA0zL+7ojA2vywHV+942WPNibPbHXd
mJSbRKCEmexySNyxAAtt267QHTyiM1kx0UB9RsD6PYOd17S6AWT1gE3nh84/YYqe88gScVai2kHg
+xNtvUb2iApKy8/nyBpVrSa7tQOSlDs0hk3ctqREA/KcUb0r2l5R3j5KJQP2iDzWGBZFb/EWyKd+
7AQiYW3WIYFVotAY+tRJLlKpmjJDWjOtz5tkDjy7mJPPsjdeIHZjFcn2UpjMVIWvuxcymOxrv0El
AttT/wDDw5BbadN4wZGKqHfpB2n6sizygb2/GIcpiJK4vbqFcGcaJLvoz4vEwG27DDt79+ZUKz37
VnkGmFt5TPAc+MQlL40aN3HbrrP+SLBGMgEL4fUbI2I/1q3SPAMuzqJFClVtuxXSAK7WwzTVQBdI
GESAvIsBRsGKwy0hPI0WHkl8JYZhjf2G3ZFEhAFErS6/6fcS+9tmn9jqJ0g7y82KSr1Bk2Oz4GVT
Hb/1pYe+myq0Mby8AWtObAkUWu9j/Quf1+ZL1GnjTh8GzST6Vd8eRM5dQUEciTvTrPmDiv8qsS/O
zvbsdSc91dmljkBvoCavWihdt4fGthGYL5SiYFJ7m1t+jPzXpi4D/eJ9gEaH7rnA9XeTsgs/Og4Y
miflZIlVX/Fw6k7aQoFUkVjG2TOD2fndf7jLxCA6ScRxSnWunIrjpuVbmpghIGC36qQ5GiS/XcAu
L5eTPHLG/+S9BRlM3GnyNAtM1iBZ5LMrZ+8UnfwBUKZXXFjAYzo6l4f1LqFM/4Y75/BlSVbq0KzT
0WgHEdOpuHW6GML+Sd0dPDK7c973WHst5mG6JBg5ohXZoxdlhl6nrhEANBNyhpvLLsPGR6+cwPor
RTMDRVuXohxY81El/D9VG6ZAJGzS7NFX7DcJAhNNSVeH5O/+37dM9lXIYMQE0KvUOWeEwXRfRJGM
ajWpk3rJF88EjeHoj2s1kuId0e+fdTvCeW9dVeNwluJ/hxfVv59Qd/TO0DlRep8QaaOkfoadUPDP
Spgc8ALsbJwZ/pQ7m5NQJ8uxwr/YN5d+EoyB/6di/rV/5mFW2mSoEjOmp4WGT7M3ei3bUpkjrUJh
Gqrp8dPKqGOuxHcKelF9s5XYLVQPXN/OHV8pGprfYRwsSnCvn9ezgI9Rplj/OoGgRMuKfEwj5uHu
/K27eoYHQ63UVGClxmOUdn7c2lyP8nBJ+0IEctduJXANk6zoXvm6cAWp/L8DCCxOo6i6vwng543h
yaeYjyFSHeYe7xEglB1X4hmv/3h1cxpDD8dK1HSGf8FuF/fAO5ycmU6jrXV2qjdW20Ou4+KIhBdl
emUfLWsPp2W0ItdD5iwN85XdQGOxf/5DpJ4FykV/CPdPOJ/9CrK55WvEtQeerFAYjh6qW9TzQOEB
PMrDZiq9mouVzj6JAQljIFMpoB5ExjpUBI+ftfUtS+S6bAeMUFTLBEQhB+D2uO7Gwz/eiN9Li5dQ
ub9WvWKIbag0A9fls0qDCn54piz6dKIHh0/EgHDYZH2kS2FW8Wfxo1YJbI7fQl0xME0EUjteSbs/
wSKvJOcm2MANsoffZUuv03QjzJE+/VtF/KS+Lbsd0kxXwMFoNFa5X9t16k2mdhqDXCYKw0SthzRR
rNOVREgVjl4EmYpjpNG6f7Q+KOKBNRzele8J33EyNc9I9MA7snh8M7gLFlz6WJuMh0HljM3qKoVW
1maTnqFotUgURey7h9jiR8aqTTo5Aosf7IWpcEGgk+r39v2TfJUT2BOSABondOv4mDU7FXHAD9DC
XLoYHLqJv1rQ0ydt/mrrLc8X6qGLtK76K9AFKyrhXrkpXsrY6BKEEEd+OUGX6W+cUBqtAA3tBm6n
/kDqOJHUjmfv+QMnwQd7JEk2Cqa8if94kOoqx4G8C0rnoSjDiivuf4km83j9rI2iCReYQZ9M3lVY
ncW4W+MyfP3MU9IMZn0um7fQ2qCbpy8ggANnWCEkpzFNZxScrHpgKggT2Z76ZNXV56EllxoRKyqN
qi5NFXCbepAmoi6mEbdpwcMY2BQTqf2BrWeJCyYuLroaDaNH18lVHYrC1TMKwXd7flZTfFgTHEbP
B1m1G0Ms/8Ey451EKYwACsHhtDxzs5zvwPzVDFSYmfrKWtHV5ISK9qc8X3C6/VZ0eX3gBIuleZ5G
jjfRJUow1ML6opaSs20vq4g1ZCIS1H+ORB+vnsGQycvf/on8yUiyWgikcmDyGAUobKhqZnPTaUIg
HEP59ivjSH5UhrQ5J7J3DOZuI/zrSs/xj/E/6WtpDIGkICJAHyf066gwW9IEMtB17FDIVkMzF/Gp
pEkZgPE25c7Tz56E5nVGHAz07xDmU5u2Xae/5yoIwIIUOgZn364fRIlLoBNmzRnB9kY4q90nvgUu
iLNh9ofphtAhZZfj1XTNMolM3Ou1gBqFLnaIJ9f5txyngD55NTZAAQS81zuLEY2Sxy+xmvcXNlwn
YjvtJCeqF+QHoqClVRxewb7OcF8uiCZarHHNe5DiPyikIBS+1LFweXIJJH6RIoaplKxCuXBf64lk
XbEqsgg0yErE7v2N5tSHjjh4LJFX/KNwS/f0yZWsYTwm2a5lUXKVrFkmYLpEekbcRVyHWBZEM4PJ
vjjKoIymEKamp0R71XmbIoLlKM5kJrXgnwwRtKsvDPdgI/VhKCa3JsXmR3S2QZ8A5w5K1qtFuHni
Ha9NNzXryCeK6NmK92aBjqh0Dt18xAcOPWgB0/H/9FiKOI9UQMI6NnJhc2+yL9kzx8WxjFK4U2hd
eL9Ls425h+tR9pQvK3zN2xDfr0OZ976SyxdvsWW5vLgs5V57mNyQNym6XtfVttvy0yBaXLfi+YSF
D3TzJepNuI3jjIRmwfYeQdo9VFsD/oUzXzRHHm+EQJ1mNE9tsVvZATCnUGsDuTDP5wH01xkJanyD
pk9XrZoclHccc5xGXHnMzaiQMuyO0/vHb2kwAhufVaUu/8bRwaOaEl3CQhu8eDK9LyU7NEmU1zVR
AzutAxcJbPO5esLogQ6Ayaxf7z7nkBVMWqOmO3l5c0fUburmrbP6h1hxEh/uAYD6NYmqdoW1wqp2
agamtgH/cyvaLhgnuBMtq3Hw9zuJAJPSM1RLJKJ38ufc5tyh6sclL/yZY47dwSzDwM70WXr3umli
jk8re9JMyq14IPKpl3uLHbdtKqM84qnzJmKeVsJDfie//t/BQtuxH/RZVxHrVs669/iC6FY+r8LZ
1ypbRRqj95zOxluAAylTtapD+OBoVoLnFQ4iBNITxOOOP9deleSWFSz+jvXYFfQYsXCMimbZcy+A
uL7LeQFZDC5+e0aLIOkMM+noTtNy03x3944luvKLmug0QYWe5Zc6BmiihcxSzOjd0wCWoFvYlHGG
ZWP9W0vjSFIe9YrHEDoAu3Bo5iBbMC8t9qb9scBeD2uHsWXJlXp+ZYqG++jKyFWQdBS+jEBlHIAS
9VK9i8frq4cDIjppl1JWfIO3Q5AxCcoN3ZT5TnM6WR60h64hHI3m3iq88synmfoyFFje++fO79ek
lJAVBuJs20bhGgUDbFF28PlOjwCaeLsErJSyO16gG1xW/K0ty2rWkIuaAvfq2Fk7xqQEIBnAV8I1
bNQrCWIbH6IcbRz+Xk3OPJKkyPioDBP5+ApeUE9NgKhMjB68fbXZKMsGAHzrFHK/ju44uinQDaey
PbgkFjT/Q+NQybs03qnFU6Fsgsx7cxswPMOE+H0HlPR3gcyoB7yld529XpF5nJgDe8cX7n/lxtpd
lW13U3UZaHoo6LyLtdRvWlLd9hPW0r+RXaMt+0i38GZw4YBGd2w4RsFaBi6ntyNY2pxgdpQXnl2G
pLKHkL8XYKJR7dJNPp55HWPfvpx30b2V0CIBs0+1MCvlVuSxgmjOEoIKZJaMRZXpu/ER4rD8YU/d
65eQr0tuEqeE3/qPMw2IFuWkVbH+NeWqMC/pXWKz2Cp5HbNZbShsBlqPBCYRrr7B1QQlEOyNWUlW
/9r/BmFY/TGUv9licXU6tNkxayXTVuGYtezqz1sT/ZBeb2XzvwdmYbQAtHOSJl8h7AmeYNAN+sRq
6p3nAmvY+jLT+UaNFuw1r7xbVQvs7G7zlcRH67BF5ZbTIywJE+y+wCGNkIc9v1ykb4iHA64RLH+T
oQbiZ5r7UTp3xqSQhWqpo8dW3+jVjMobjlxQKGHOBAcizceswTf1nb/2MHA3pgyQB6unk40EaILY
m1kmJoXtukgX9GeWmwD2tnZDQ9QLN4LmzivhMqR1MPhjkO6fTKRQKw/C0m1P9muG9nb5gw+2f+8n
p3+6KsBg1XyfXX1PGlpW9/HDedJyvrg0sQApbtzTPunXGtVBMAAR3PQ+byRD2Tf9kV9Gb8F5vAUy
YAWuJ35R8ChP6WEzuiCrCR/pne0sBfxQrrzoDtFDvD3G14IV6GCUtV+3MhqVzn2oGIQYD7lAhuC0
SNJmkS7m+FpbENhEGI54u1Xnho9u3llHoc66yLald7vcfHWMxjolCKlSi70DtedrHyqbMJqen0Nd
mWgVegQbtLeTZEgnuBQ+nMqVVj7lsBJYQQ4wMNNOfLxPRjpgvDY6IJgLYiJg8IX9Fy4dwz23kFbM
qQHnVb/YFBlFpAM2I9TU/xja4DtwMICckzZpkGXutUPKNmody9lWqU/I+zPW7hKZWnaUNUpKK2Bj
gj/TQNgK8EuJazYFGv0XT2K0d66/MHonHKAG+kqxDsMVzdtlqClB4TBEXWH3Dm3aN5zndTFRY2oo
ZujRUF+R225cyQIscM0zi71akrEwWl8uK4iKrYH9D8oTl377AM6nSGgoPs7NAYln+50rwrhshqTY
reJ4DQD0ZImSErPOF34JGAO42Pn77aabiXN0oRi3rXnRb3oxuWjubwnQuOMteQqkmqhU0Ndz03cX
ZtoVnEV5o6glQWEERt9bDuwKut7EYDZXodS4GXMa+/m2ct6oF0P/ROBLDLgRHpJEbey00sH2yEGH
23Hy+TrJim41BvJ2Xje0Qnb2jy4ciQ919kMhd5jGSyrLwQ1Ju6S8rH702jibUrCCAsffdzBkfMJ4
BtpWy1XBXBdt2LBkqKKEmTkKorAex3YzN7mTUxXg4TBgphVlp/+P61hDfyjNrolcQ2MzcwH6Z1Uu
iI4FecPxlI6prWxvAKNfIlbTakBdcLiIkdvwMwKq2OQo0KRdFjzJCJLtZ1c2oWt1Llqvc1P1TWAZ
uEt2yTA3YOnpcUDobguWGy+OLZTDPMlyRyM10o95Sv+rBbG8/Bx1iFVeT2ia9yZGFRUpIYqDrx2k
kY96Nzg6y34zLkq370PfNsVWOt4zrQ9N59w5wmaS6c0ysvnHmJUw27cPYLEOYmlE3PRF0RpP+pqC
RDD/wfuLW5FU+EY6sIHyLrMIryZDlh6sgMmkf1UJyhJ5utcjy5/FcOc90hLL8p/3bcnDmg72awK/
Oj+RlyUzFFRVhVFYY2nEE8p69831CvHiGDDj+XZsGFg3+8eY5RtyNc6cyjWPpu0z2pq7fVz06Y76
su7DSV2R5Sjd6VHSfhM1Qz2LHUKurYTZCG7QAI43+Xak1JL5EG4UKnR2UwDI1ktigzpVkjkUF6U8
WYqGq3QVNA7T2vvcMAlIvp0yxxvoEx/oh+sLOza9raTKEN22NeTzEgsWpO5GZFdCYRKbeCiCkC+e
sMKEDfhbtpARWsRtyRugOgAyiCK4D1sJXZ+UqYQ+k2YAgzDgzJa4Z95V3P7xE6u1hbDOkSDOHaar
Xuia73jiptbqRsvu6kbGRdERAdFtZXoDWQr/8rRTA0ykcsTGIJaxqy2+Bx19Ijkn7hhJ0o5EaMvl
wUnjcgP/Pl4Y+F4kTw2Otn45qxpGJH4/knPziK8aDfv0zIfL3lnSYnbMd0kFWEwPz9M6+MaTWzSm
chK0CijtyaNOkDuQd+UkFzC5ZHN1HlRS2iu9oXvkbVQHf7uMDwLxPspW8yMy1rh5C3RCLQ/ve4ia
wuA99uLiTeR24TmgHDnkU/IFOqHMtndE/5WdUa8hFaIPOir1OfE3I6hIQ8yamUYY0SpscvqNH3Nd
RG0DP5lF1HwyOPYU5kKAboZ1UtkAKPVZRTIGpMNp+Ogxws/RAR/RiwNi1uRKOalpzx1ZTW1qnxae
kJMv6jxYK9v4STMWbhPZylEMP+nZ5mPNghRjjL10xt8HnNEjWL0LtzBgBPO81Y3bpx2f9bjdQkRj
N9KAaxo0fB/RHfHLqgHYSUhikRKRqkq0vGxQRCw4SLFRQoFwUuRabiu9Zxm7np85lb5M6+LjAl9E
e7S+MS1dHz/KUuaTdtsrA0J88o6IQmt1eWNDRzda1ioDbCHH1WS+jq/c2MU7IcExVGRbLIm7CwX6
hU1vkCmqTQFFF9UybwImhXf0+zBLIdflA/1yIgxRGf3UDwAwojrUfZwQ9ABzRruWSo0hEUtKn6AQ
n4vmUJuBat5208B5JKH0cJqqsAzJdr4seMp4XPpGIUwcM/ppwDKvY5kV4mdyKcUcG/lG81fFSVfB
EQHPRybdPsbDOCcL4yFyb/L/eqTbxvR12+Xqa/qmwl4AftzKGWT8SBwnFeuCmcutUVGCqo8nOAyR
C5gIjGIRr/ta/t9tno2eFIRDfWbChPAFAtZ/9euKuaErgztqhFaycELxpuk3A3jkMo7OkxfDreqQ
zURGfJj0e1mlpW/V2JHy8dWz6tKrddbQYk/pcCx900WPe7HTjfBhQWQkoiyQltWDTEfeFrEkZKFD
6YV7cbx1rOfFV8jnz07l5H+e3+J60YsrnMwoIxY7Gm/JbA24y5ZF+PrL113uX2xcfxiPiCnJxtLS
blkmZblEnUIOjqCe8dAXdaiBsH0KECtFhNPwafQGZXQY4UBA0FIOZRtClobyIz0xn9R7nBn5ORUv
Us2kRzJfq19aC3bgnE0V1KrnciLWXB/+pT/PB65rSfAfacudRWn1UmyfaoNrISHIM0iyYP6UbsWo
CRfj6pTdSDlD/QNMRRvfvCqXQxCjmDclGcvj8lep6zy4OOq42gJ1BnwzUoxyo2Ssysi0EB/Tdnkk
bNBCbNOeC5P8nRAEniCQjQRtRzrsgNRKWebQSW4TA7Xcg/kcVTcsevGomHNBsEUWvpeQvJdQrcZ8
lNSKZzUwa9mEPdo4HY7uk9WEo+sxajf01w/RqijGRMp9vnpmQdiyLr4Q2AwBhSLUPSYcUTg1qRbW
jFFpxlodNxuw6jMrAqeJ3c09UiAuAMVafEQsc7LW1pPdiV4EOd0Bitc+G6EJQhMLqt+DCnTYd45e
qGD5OnLhB5G5sqfWb4pp59t7MsPzlKSQOhje42EY8rFF6sK6j9m3qX5OJSJ5rE+c9TNHw4rROuNX
YTpyKuAIFknbIYqU6mXusPXLWUxgy1wuJbbR0wFVZG7gSUXwk6KN+iTsCZ4SzSXRolsIWZ0WbCNl
GRO3sLLa3h/PIySPMuCYANZFkYFFj6V5Ipx9oOwiM1CsPUag8iTr1nW3aneZUuyPLw0smar5qDIX
W615bFoFenweam4WzwgfosdtewhMBr74xzdqzeea4LxeZKpRP+6+lEH4/veAONAJ1BvcRwQ0Bw1Z
x0LiT+D2wI9064YbStBQZ4IHr1PzKOSUnD43qCkv3Usza2nODwGVcttx6rpad9ET+eW/JnHIjnlj
xEmuyraLhKc18v1VaJHpSIbk5r9I31C5RwXZ94SSZMO1pqb/51eP94e0O9mKwodEnc34lMtvgHO+
aFEv0D4OZkuSgIdKtWHwAItG3NyBrWtpjv0WqykqXxTM18Kw2WQeeuF3/yGqmDkTlandDP/tHhzK
bzZsxgRrzqS7qxozbuzX55xnPEMcFge4QISEGo6LGKDxIdjuiuC4kzAt75ZyuMB/w7yN72avHsNv
LdSy4dVYjI8gM0olw/npli/0LwlqtGXT6ywYa20REpFIl6+1Bw37QheLIdL6zjwIZzlReaHHZzVt
MDmJZ1/yg1VyoepFshkw+OXK1orCvjpKPP+XCLIf/dNY7FY+6YjqKv8eQe19UZGcSRWUQ8t6CNiv
5TXUN4O86f6RIYgilkONfzcHumNhAjaUG4SC7YhJ9i1gT2aT4+LEf9nUQr7zNskEUzbq2r6Lbgw1
Vu4/b1y3AxxqnMfqnQRKeOv40sPNWA4/SzpSlF8fwGyaFpM07vebLkCMzKxHQ0QP4SPijOtCA3dD
SADgR/4PRgboTjrwVFv/ukQWVGb5zaH/NR5rVR8I5Dz2lIv1uFBbJJku2APYRUlRMPGF9a1ofRzL
5DDbDxYFFQqVIWzbO4rF4JCnWeNLWlxLibvZtgV2rXmuEPODK61oj6tiXl1H1w3Pmb+twobYzpYQ
RQGvkvjRBz9EHRTUnaHVGzSsGIcNbDj5+RkrRMpGKPAzWri+vP4SAgLdpI5IHUwFqGC680BIbIyI
zbwnQuHYFyXwcsBWoT/6c2PnwnygHr1weLlWzraH/KJPOAQajfMzNHjYpJ4NUEMDpj/DoyGqyGtb
OScOgV9TnTT3wAkA+j32lP7DbCycqETcTfFBhswEHaRTWfzLGowmvFjUWMPpd1GlexUluMaNMqMJ
luwJkAuSj0Ty4xUkQ5KuOQRP6U98g3YORQX6vZoBE6tmyCgJzlcViaO0okKZB4kEqHsozADaIY4E
Jxu6gl82BpP/w4mgwyO+tnO1nwbOrczYUjdXp8xlhgEpQN6/6bxk+urzJ0uJmDH2OArEa5d8tGMr
GGyA0zuyRDYe+ww1vYPaisF8rdXdF4YRNJUzTvOdmy8+rdSZdPxVlai6LyhUzla9U+cvBrVLYsHQ
ipruBGZ83zVLWVVKYmKIoJpMHqnIF4F5XZmgscvbSwofST4quIDF0i/QI5rhB0R9ciOLwW+xH4lM
gFzGNTtUlrMepI7z5eK506PuKSYSagMX5oDTNqBOHTndnji6Go7J+ON22HelFKfcrt9KokDSeElb
NUyQJmRP7qhG38SlUqX/hzoyfOpbEPyub9F1sMei7PaDaeeTL+y822PF8t6Ro2eDNpAIa0jJhOnK
ZF4ruRFMGJ+APQlG0A8hxwLWsSKEtkUXdcWyAiz6Cxd/foKVrAS37SfjVxKLXCWkK2sjxkK5H20B
12jRC1Wxr5bIeeAEMDyAIYqCLFxGC7A6DyK8As9gCXiVRQn+o1Qw3yYPpX5HbfA8+qp/JZw/jRWA
xuwreyYh9u1cXDFCeE0SMhFp98GUmyiY8uqByalxN/YeyXgfElf120MiQnI5PFLuV0+aLvtNW2Ld
wMkvER2RTij5ivjMRyxFHcT0bXolPa2tXpzIbRVPG4PJ8i7xeJNMdd4gNQWwkTzQ6ogeOLU9MbdO
zaDeTt9DoS1iOkJS48z9ho5VdehoV8xr0sKG0TsakaLI8MoFyOzrQDOCKIVpObPqNNwzOWoSRB77
EfHmp7kiaQjcQ2oK723dKkNLrGvi7acq/102Z6Q2Jrtr8ABqW2XM221GkKHhnUV+OWau/X0iyCwp
LYkmCpdGd+3iWk9PaYcFHSGoopm8kfCbEnpIjlQ6UcwsD752fXTsnlRIlBa7QrA/SBUA//6i9esl
pLCrRjFTwuVBY4a6MT+VHtFDp3RsAyxiAg4O+fCb7HnkVWDPd5BEx8YLrLD4UNANA7dzzSxtllGW
yDltbYJQbGHhZDnuKXdP+3cRssF94EnHg8a160F8Gbvxi2VEPfiYx7yAp6tKdf0GiBm2EV7vcgpM
87aVwv3cVyDIRx04s8OSSrJq0lIXTUFrKpAQxDmtOkIo9fBSQMdyvsbIzXsQPW7hRJ3EkynWIJAZ
Odjn1QmT04yQygP2c6eZ2K702hYVXu+WCh0UOAPxS6pMh/5SXUIf4nTYpOlaN4uVbfhTL+FeJgsC
o7urSZ/jZsTpTCzS6D+sqRjU21JxBkn0tberkFZkMWYMKFY88Ihm/6gTVKbbjViqV7oWMpgsUO8q
L8STGofSeE05pxEOn48SySWC7v77TP4Sr+reWxHLGajFg6dRpfkUdGfdQ7pSpIlpBjbe/PkK2rCI
uRKcOerJHO1d+O9z/WVmankELcmbqg57zavjYcy3GBDNZN+WfRvKCzGnH7+YW9J3KZcu4nvlC6XV
j1P6fLNKtYpQT3p1RtpyoD+Ah8AWakHwsKIbzOuwsnpmOspuJkYNIMNdlZuXFaOLpjls1/4TPrRa
z1xfbab12ZePRY5ZdPycM83cjEkCBRwcRVqhjStk3ZzdMEHHYb54Vf5UZdleU+jfPV6KJ/hY1zdE
ze6pM+uZjzcLYMhiM5B8fuU+EOK1VQ7rimmzH5CadSeKyawOkogjYljBhcnkhSk8uNldBOBnjSma
thZmnhW09+TkQ7FeSmlk6HBvha0LoOa6dj1tQr5ReYHruuPqfb7N93HckfqAydX04cMo3GXcnm2h
qzFnF047YxmOqhwDxpGlJgAEOoKyglSDosqgwX6k4U4QFYAf2MaR/BkhrC91pOy9NAIe9HWvkRGt
zVhRw38ZGSJKMd7Y+UvvpjDModTJbXJ2NIBjlytVdMeW3MA+GDajGV0Fq+bTcAKYTirWeNNVNnQr
m5BFvV/qHio0dWvBWlBoh84CmHD0/6cmUf7mlFshVlZV5KR7BewN2qrC75d9WMwiYMqSHmtJuM4R
2KzU18UWlLvkPaG6vGbUI3mHCLberfaS3Btra97JgwV64VXuIzk0OdFqZDlyWxgfepMVO1gXGh0b
enSFT734h4f3Y4deUk2CUf1R98v4JKTD3uXcPgtc4y4VkeMYZyOS4CtoRK67QktnimLRFFTMnyxw
SL7fhP42f84GeI99YIuJ1LlOyd/Ay3HGjDdpek8xW+BwXdOHqyR6kR7pkyIRNVuaHepe6k5U1w1y
JYYa8N0Fx11l0MSw/gxZdPFctwEwyCF6285+zkbHtycQuFo4QQZuT2VXHxVSYhDugmtHcrxjMPcB
LDxVkXgACW04r4ecalvrP/jxgVtKKbqilTL2wJV5rGsFX2ZXGXjTqWn5C7CIJZzA0Kbq7lHPKl0+
wPhlVevt67yTaKe2lAf7yRUUl7sR9WdGlttQ4BwqwT/uYw3wZqRncKusxqekMj1PPGlsesW51qYg
lUvCmhoI999wy18YEmBWDDdWqAhYOmK0Zk+AUL+13Iq3tKLBMRTRCsYFtOaRuGIvVOFOpSJlFJxC
Ljwt0hLeK8EdO41/YOVhf1kJnSonh5z9bLFQqXKm1xVai6moGwVq53AeMr7zL0iuGRYclBiX4U3x
2hfUM1CeJYmzjDHO5lgabbeGmvG21M5qEq5x/TFtgcd/gSd7m/xkCnQdoA7CHYgEP4U9WWh4ir1B
QYP87vCxmUmmzDY5yWgk/kxJLyxq732DO6ryjUTTfPwocTTcDwPHthxfHR9ywrz+nUi1oO61VNlb
p9N86FVVPfhywKampfcPOjBWNnJBolXA5mUQcTKOvBBGEGRTwp2fO/6HmWzIW6v8WhwSCgS4CtHo
wjYaYqQV/yFOR0T3oWCb0qJJbM4S8HTqQ/d07MxhFPIb/Q8ZcBF4Aoakf6UoNj7ggTkTK/iYnWSv
3U5QPZ9Pymq3WzM/hglgIHnzD5WkOSR4Ym/fVoCB4kTVc1RFtgTXktiaV7d6vt6alJkNIv7V0aKu
cWCdKx8okXJnxDv9fGSmcvho0B6pR2u6D7q+k/1UgsAdlbx5wHlVpSVJPn+Fm+uplyrCqa/BYi5F
ZtSXlhN0rdtwpVOW5mxBopWJIkxK/L7PYLsLZr26ykAO7o4nqbSZnJtFACdmPwVpnKnS6PKNuFV9
c3oFWfjvlBLcrALM6hCmoPOI4gCK/boON59EtVYZVEoDVGQFVaNfWXV3dlXN0eSaR5PE1BIeZ3Qb
VsEzfl21+Uil+5HS5px594wDaVuOj9/Z6eR3dxkvMAszqSW0qNam0RQqZ9rzCYoUI5t5K0pPxQ/7
S/dvfYpsUbkK/AZuqqPP65yFpuhAuekzh8g8s6R+pBKO9KQNnvl6I++0gp/TX3DYMRLnp0FUcYPb
hSjW8Es/yQ/F/jigfJiuGvkyIkQ7fBhkTgoVnei4/ASWPwxwW0m+1hH4EM8D9akIBfo/FWQgXILH
4UamzvKuevbrZqhg7pJnI0ywMaO+2oLzW6lmbnB5/gfKv9/yJAwR8ic/rKy2BIM7fGviZsColmsk
xEcV3qa4HkI5g5IEBgPmA/1FHWGuOFKFy4aJpOeeUJ/k3QZy/AUVq4KaqzsE7KiKjoGRvlYtxAXv
PkmmDj+Un44X8GqkIO7srlWetKeVbWAlffL5AwQBLxS5JxrsAJ+PCSwNeqdojAbuDOEqFL0aQrx3
Ly9RIekBbIIKJZILlJPI7lGZxOTW3QZE+3venM74wYUzsjQzVEVhTw5r00X3bxQVJhj8DDhDjO47
qfgNo4x4nW8jgX7fNc6FwbsWbMBe6GrNgzyPihfTxOtyNw/RIEHzqiv6odQZcpsg1EwT/xAXYtol
7XJrny3X2rnIiLwC1Ay7UqdOvJX5Y6vwSopxaC9ASt6aYOHgdsesFkIg3/7OkDG8jAhP/RpmFrsS
WADucpERasI8HociMyGkKqT4PNo+nrHm5xZhu61q5lpo1EIwB2hoGhIOOH2Z7sbeXzCV2PDBBuI7
NANdqOwc3x21taZp564lGFu33msIhXu47S8w2RIiNavo3OzI1CsaLJdB0za1gBxOUWESqRXRKQOp
wMfiJf/xHw79vTbKyVI+0vmvwIFPCGe+Kel0PthKlzCl+2laVfb8breJIxLobYKMFtyy+tEporRu
oLEfTXPNDmsYB6LehJQspPcmpRefD+asl5lWKgHhfqK/WkBj3rEFaRRi8XA3/CkoSvyG4Y1el2lq
kFxDagPFpwFUZCdEneuMNRKGzEoMP0k51P1t8ZByWiDTO6t8WOilQMhBj+cvgCGbahyFUyk6Qfsk
HIT4GOa9qRKoHVh9OQSiAyPiutakWxv1XuS1akxcO0upbqWXzfAYQONCqLj4bnv6m1rmOIvHLWZN
sTDcoY55NH++FUOtpPdGombYavQljWssqbGxV6Q957uzc9MHfW0N2ngZoVu/0bsVsFA6jnJvp56f
MzRJhQGK0d0vJm7vqDY635cdAwasUQpOz8C1WntYnlcTcV4eoqjDQ9C6Tdl00YKceE6T500MAuct
JuQjCceU46cQyrQB2t55ngwH7iIYiv5s+dgZIpRBAsDOZ1VPn4btzdwCss7hithoPaHotG7J5FBx
k2TkEbvm/9u5UMp0lqAHlq0dO4UNvcTd7cFOKzIal5W9Uy7zkG+fmjVYjfioUunNAY6KWUIiwXUP
2Zfy/HBy60Adm5aeEynwrxw7CAr8QuuN3fuf1AID/dA9isajsaThSonLeGHzERMpuymF2AUZ+mJC
Oz6bVNl98SW40vgKssGSZ2BJ4fBkgJAUwjKhTKPEO304ZNu5Iqv7xTuNhPLgf2ljaNq37zRY5Myk
l2kLWRl0PWJC/H7Xsg9AHxZbafbba6os2rQ50U0D+NWkk1CSG4w5xdggSM35UMWm71VHKunJZFLZ
F/TfsCxS93McyGu0KIJzaddv1DJ7x9sYwTat9sb0775tgN1as73RmLFE8G0NG4+P341gcdMv0bBp
jpn2y5L5o8FcYV9T9hNc4S12PH2YpR/h+ER80wZ12LpDPMw7IlPh1EnMUnZYazcAVCaouTlCZmNU
GTLWVfAVM9wKBXoH2Q9DDswtxkkcn67zDgQSSqQPGKC9pHpCjpeumPJXyQZhSAI7H6TwjwcH2ZQ4
cyn3/yc0K6+zqZ32e/tY7FXHkdCGv8VutM1WU+eZ9tX03mWAhX5CUu47rLAnjwYZCtZPquXxuEJi
HbSCuPsAlgxpBwD/2nBjA/YcX6VtL9Tviam+Xs9r9v5K3vFfkHMvN6wXm/ZM4zWfYbyZ40LJDGnM
mA2dCUeBwBwth4uchNCV8/DwTPvYYZqng+oia/aQd4EqeggpcjnGcoAZBOlOknFZ4RaxHbSCmB+v
/k+IlW2EABwSW55ZKPJjzfbnQojIZz5yt3RdXg/RghY4afIq8Ji4WsWY/loy3XVfvAjDrbs5VBHJ
ltETXuo2R3dAxJcMy7QIy7wCJuQAJqmsEWg7mLJV3eMwrlQgejqJHP4Kv2qF50cRz7DST6sYX3HX
RHJm1sNFRToT3jr4mB+a0Lc4+ETnQrxUjYqf9kVIiHmlrbZ/+ioA95GSIIYvNfMlPUie+YwU1tck
WXw/aV+jJSQAVGDCgGtnM4JG0SU9XhA3cGwL5dwSP00oEJnm5tVDMUkPEcU/nAvaiV40B63TbXiO
n6JVa65i5NPON5MOKb9Sw0V78t7Edd3mx3OiMdPbj5iUu4VQ5hKdA5TvWIjAzypyi8H43Md9oRhL
a35+QC5eeTXhRywYmbCKbmE52wurSgrqxZNCm698qaxXmU9T0wz4JMQ5/aIuTkeAosSN+pmpEQ8j
OHNfIGonFRL88S4KGPg8V/Cah2HT/yBWwYYRE/cWM+NecmOJLqPSRc0oV6wy/+6z5rtm+q1C11Wd
hAgZ9ajyn0fhYTu1XUm1JM/VBKsBwnZur81jw8ilYiEcQ1oY4ihxUMMNw8Ln2zRvUZzj+/+1kKuj
7gk08HxpdyqLxMRHl4pS/i1pVhFqu7pN2vcB+ZRh9vV057hn67c+49oFIbOeU1RDh/Xsg1aJXZ73
yD6HjABVCthM9MaMOuataowSCankT/UnPKvVBmrVFkaHnymmMiDBgHtNhkhzNOo91zJJrOotKwJo
kID3PdnBLUt9rPAM3iVCTscVmww5JVbGNYTY+4HJ9RZ7oPb6MveK6WyLOJd2X1J/kMDppxqpP5m3
NX+Aq2F4De36wvP/g1FrDm6tB9O7e095FIvt4+l7PRZP7vt6BBxe4s7AAJJXl1l0mVsxPMRXRq3o
7sRVW2tnHKzUszQ1eqF1/VEasD48oHWiDnTNNRUz94aUTP9MvV1DHb7mY297698EEde4xvmgdojH
iBk2rHniY/xoysP+7w5oRc24Q7HQ4a6MR2vyQRvoqZkWbcH2IdpJxWcBsdrC4lVPmK1jkj1aYUQn
4I+vjyejeQtjzsFpE3gQR+qTwrX8ckzCEJxfMrKWOygcCkoKkaitLcx1p068wMCYxo+PqcGwBQrD
0mHq/5bmx3HzqDTXkBQXgIWNEO6fP78yaWy+Sm/NP+rGgZxE36kGpobDd2XTwrljS+LUmHBG92Nt
OPT7knIX0hTpGyNvyzhJ/6YXXhEyqaYEDs3pkWxvJz+NOdKdAlAHNHWAo06jqfI/++FgysjLm7VV
HWjvwdjYWGYKpcJbgLYivBK+Edqmxxx7uYrJ2kpwlymPrjuVxvguTmZAaY4TrudtG9s6Rre9XLdL
5Ycz2SQs1BXzmxjP97ThDzbObXpJbgRi75OyctyaGkC3WtVtYiFZPi7kV2Xk04VyqDxkH+8JRR48
Wilj2TqtOSdKNfTSaMlavcR9E1YUhfs4Jo5opo1cLAZDB7RAFBTKABFMUG9znpFF7DVRlkZryyHy
CULKMALOG0S8Rg+O5P6WJbDYrxctU3IhHshjsBfXzywBrGYpXO90Oo70cQxijGIUdb8+ASBrQeNB
4ZIi4GobmFlxEw5k+ckKbgaUpI6PPMpNOd6SP8JNhVas5u4SfkinmNjX0is3VucvGF6dxRJOdFR4
4trN0T/r+Uf4PZ1WNlelcYKkvPJdAcxuqKDdlIMDtUf2pRGDarCRBD/IQmzY+4gFJVgsfEHOUtAr
CDh29PhWn3YZigcq7qt9gXygY3ZuwDFkF9CgqqlyXi5XCesPmzgSjAVauMxD1Tu/aaZLlOry5OhI
+DZRSajiOuVoMmN3N8Pg/buEOs3f2XtpFNMMhQ7UvJDHjwPKFxdh7RaTdhZBMSOQ7az9FpkUz18Z
JYQTie4ufEVvVv0yCbdt6TNeKWx1U6LGK2FDLjgcOlHjo75Jfp+W/rWTpNsX7QQFTE5bz/jAwcm+
3r0B5H47tOTQBhlqzdxLfagQiTLm8RJXhOtP+v6jSoWyljfx5JZ+r7FPBq5WpgB5IFR4a2lCTNc5
B7nsApRRsDhfriqiQ9txA+068L0htWbtwNUFj8iBqklLq1/qZ5T7uuelrtkJM/Lr9GFPXPXgHaDR
wO4K89N2Oiav9SH+jIYm/PrEhGCJq8468kl6/nwx8W2zgPdR+ZkkJq1mHCCJj/WkXz44QlgIPcVK
0iJO0HSIjHpeTrad6LHspFqWFtw/DXuZ/Ude4Hl97fOa074fDpOvFVbIwqipIWPir22tu32DK4jF
fwmtQ/bTiyUTtAk8P+4ea+p120iceksPugtyUU+x1qhn7ezgbfqmmMw1tvAnOHXtifuyAlEUh9Al
ODRPPWRY+yhXztaF4xCV0FHBqa9tAVChI5K4ZmecURlA5b3erM7S5araA/hgrxSZTraqAwoKEmy5
C+OOIT5p8Ujs/No4T0/PujTObKED3R7y6gSXGeWDKBiUs/cJG/wJJXwL3z8gPSoQwzltf4ofHHE4
idbn233N2U+OJujqBZ2zQdDqHX3Xck9P+CtAc2mygGbqh4+eyIyFjnChm2scUwyshXxDV5vHZgPv
5UoPBhUn8QmM4M1oCfchoklUYQ7WeFrApuuPYQzp2PZLaNSVe6zFWaNw4jsiC5YYcCx51PfjZxY9
dmHXL+mt0L5W+Tf27JRceHfwO+A2w9k4sGk6ZtOWZ1xExTqpOL7D1uWJKrBrzfAhTSjTAqkSK9Ym
7mNCwSOHz0exzLwrJWIicuvyLzFbfUyKyWNeAY1qC36j7iofXCuRddUePMUdwHK9fkxA/Io1blP0
dubcLuPpMQaR6Eyi0D7P126RCTA1m7CRVaCCv8dcP2XPq0vJb9bCdTDc1KZYD8Xx3+fbPZq1+Fsz
z07tyACZLSjMoB/4v65DeqvjpBaxJaLW8aOVgD+PjbP3EfAru+egf6kZddzf5vY7xRJ+BHD662GX
tmK5wvhWcSCEzmr5Hx5Rift9moOydU/jj5q+OCIc+e0x/gwJl5vYuJU1by6oci3fDaq2NevzbXul
WPud7dcbDX1yy4STmHfyHtDk0rU/fNllY1zEmvFs2eEqo5PLcbGw7eoy6W15JWVJHMO4nx32gYHU
U88/pdqXuBxrk1NFd5kUgf6AXf1zEEUHgTb368+MywGE0utkMLM7gFUFYjF2HbzZx/1gu/268hW8
pGwj6999yWBKZU6qphgzJI/AptRZVD/Pnr8bOYJGv/xywRqF3Xy1N1aRaf8ndrPhhDhsYDBYQ3Cf
HIgLjT/YKXDn6yULOEmw+aLE/vaonsrc+heqDT2dwR8U9S10bhB9J+Wd0hu5m0yUFPMqUIErlgqi
GJ5j9uZUO8xP16oQZb5kPXb0PM3issRn/6ixQcek6Iuxh5vc/q4yDVmeghG89AF4blO5Pv1E8bfW
WyBGtswLVzgwiXH024+vk8zxCpGhZW08qYeQO6d9xxYgGdmQ8wJsf1Me0D/jZCUdWOTOVkWrHhMI
2PFAEc6OJGsdMPh5HLwFGgYPHUhg+LkMMIvDcMWcJO5G1gQ3eZxOid4+8d9Q3hc9Bj7+0miO+Gwq
tKif9p/Vk8Nhxz8/jzsNxKonAozX/dgj0cuC8nQYqZGMnbQi8Vv/vnK2XxcUWPc9lEqmyV+2G0wo
7SyOaCY/k7khx0Zz2iZqJGIjl35BRtiwLaNWzWkdqK4Xu1f7TFIaazcEkdrg+PcYrCSS+SeJua0l
6EdlsPU/Yv3K73nANCC0VpOusOhxYkPQspsgWhkCOSiS7X8acUTxRB+flrYXXL+MVq5f2DDpqvKA
ZaArJU1t4LjUZDLnOjz0XB8MZZAxqB+kCo/yo2AFjRB3SOaBEM/ROG+i7rFpvaJ8Pu/PGvMbjEfZ
73A95fdpV6sDl58K8kkYAuq5bQDjVAU94c0zdTLck9GUEc3aQ5sJyPUP3Jet/nEiIb80u2BTf/Yo
B8Pih+olPkgogUAaJKl+dXKn53aOFjTBgo5iredThJZ9DH1LEWUTx0sH/hKgDuZYpduW/e0HiROF
QfT5+RLQsSkEl7/lyfYTboY0L77l9S9Y6RTwrGc0BekHb8GgEMzW2o9agQLjrs4mBHMvuhgvGXdm
X5fmy35VQF+ftGw4EeIjfmoxp64GgP+kVJ3PdIgkNI2xs7dfZeQTQH5JT0egEe82VzR1pUjA/VEC
ja1AdAZB/W7UYVgQzzpuvW7Dh6bx72afaXEWB4w4LkG5q4Dy8n0a5dkLmDxfXMTjQjr+bsk7+wYR
ZRgjncahtJAcsdj1A9JrBEauE5IhZUA1PHutL95GaxxCeM13AIK37dkutHoShLDaQU+sIqifoz8s
B/huajWeZs1K+xplt/+jWKmsfseTDUnE7Uwd7p8IGMnqJMZNeyZaR+GdeevtNZ4WoXMlfUTtdzLp
xOKwkgeR8biOSxYUlJeRBvmyKWHnbFiNgqPTG4K1tcj1kXja5O2LcMWrqMZp/9uwynPZA+Vc1RXl
qjsEKPemlF+Ww2aoMZIc97ykyIWYvSFcnc6IjTwLxMHwANH/18J4llm4Rd+tYnuv6zAOwmWAfGMu
RciqRuRvZM2nyjIWHzCnkXavDRUbeDtn2WHUuZNYwHeqlr+sdaDJkW65SvKEy5119LbiX3ibQcpH
XLzmC1YBkswbLtk9zIoRysdToOYjkwWqF5SvxEj4z7aAVCjM4wfMFf3wqXmAfc5mKsHHBVHymAbK
Q9eXPIPlUrLidqbjbO6HjuzWXzBHgf0o62eSRS7slO2QqwGHF3GzTla4+i6QK1ZIMPM9QqUKixBA
oVL+rW9cRrBpgODITwTmISW3pV5CsLHfzAmw+LBGtNRuX3qoKpWU6Y3WNFM3QxyZ0gY2TsRALrD+
pctdhoeUOWUGyrkSnSAoyLCkkrNKIBfN0ipHRkGNR9yTw0cyPrFnBd46ODl3npUeM/mq11O3PRs+
KG/nNoZzRT9zaR8/GtdvBvbxWy0783HA/eBTTe2i1VU56xo58BTv78fZc+Z8XFbbyhJRaKo/HNpT
dulJdvUH+WHUIjqGqR1TbnVTRJ+3xyPwNwd1was8kCyK8Gc4Wg2JN2AQhrbjMcpZE77+DlHUaVxO
BVVcWcN48ZA2ybOm83Cr+8xK0dULCYt0UJIjmAQlriXA5VLTAvEi5jPLH3p8Sjy7ja2AjQhr8/R/
3rrQeg4xBiKNPioNKqf6jdfTvz5pCmeYVljSiVMJPBLrsk5sT3bBUqjOp6f8WVaqWpO4PiQ2NMqL
rEN4X0Ti/YbPxjoSQgS553X8Vtqmb96eCBXEyu8ZFToBbtZ6EsJ+yN8QrsKN20uB0Z1C7vXedBrC
abJMIyyUNtYiVBAJ5PwmKpMxky/GoB0r7HGYhVxbwRS8f7MiNDoUX457LRAZW7P93SnXLIA0ksbB
iCRWVWhCvJq5wMYQ+7Zlsh+7s/uiDX0G4oKPf7bslM8YBPpceqPDX14DdS+9NfHfi8BYIggOP4WC
AsXdWYofPSnNHvzOdncECC8cjlHnkCVu4+cOzy/cXSiFk1cjyLkgIEtpl1BieSW5fq68GxgajkCu
+bEj9wSn+JHIFmH2g7MSHy1etJi1afeM5GvElOP70ERs6EA0pTrmfnSFHEZ3O7E/4z3sEjjpDU0w
UfTzZrbnynlOx3NGgDeKkuNYvFM5NyXQnRsv685PWCiRYxqCoj1BeLvceJ3jldqQjOeD+mAZn0Hy
M7KzbXsfDGX+4T7Wpohs1+7/vDi0Vylh94bVEolCXslqrNkeilEv85PQcTY8kdtA83up+awA9Pun
YVpdvvJWUCFTa6KMcs6C64s8xZARImOkKuuv5hNDW74BgJ2FIVA0gd0ZRGlPDoXgCttCJxpsaich
MWns8LVpDYbzFuppOCHpwHVkEumB8JE4Gxa1PdDUHxO+3KJhFzyjdior2ZSH4ZQGkYDyuzQIySqZ
SHTrAuhYqIrfKqXzdI1IyHQRn5LzIw7027xT4fJplaRyHzKWoAqOIoytssykPpYJuTF6JCM5cGX5
iJzmaVjxAIUVYO6f7F1DVUQUYz6U0x/y1Lr/kKIy0ktbY02cOmHC4K4kLbs0F4JmSy/w1FGXCp89
ktoM8Ome+s29RnTnRFjKWzKynYwjEvkNU3LV1tRRvU1AL9+mgNkKhoX/t7dyO3RhENghx1XhWebj
J88P7+8FdTacF8rbQxT3vZ6P7ap3UF/9mjxhF6qyiHlayEtqtzVORvLsedK70yDaNPIMh03zwHok
x+ZgdbescIh6ZOvWAezSmXD08p9REghO1Au9M9f5g67XAsCdytrUKti3h7XQj2S71tJ0aIrm7vRn
nM4GIYCfmT+jFmiUgSmojtk8pKi8P1HA/KkBijlbhvUHwn6g5kGs0iRL2KkYHi4nfpp8vN7n2fbd
bS0qof5lbENAFBkzi0904riL7Rr8u3AMd7tkfyN4Bkhvz2fFs1flp4c+9CYaI8HIXkC4Nl05R9p3
7EsnDG1M2qmQCAaTCZl+Sx4sk+guJimU6ZpAxEUTb6tfc/qeCVmN5j4HbbSsLA/GDxsLJRJEnAEz
Pn1GrNlFrXKk2n9UGI3sTnMJuthAk0xSjsPsilq6J4XRKBhPeVoXqSQpz0UfejJBUgX5C5JtKkux
HBG2EK3riO9lvNocKisCCggchz76LA7nHBO7DmbJNlAaHOtX8L5XoA/gR/IdmCZfJWQlwtYt0pO1
eA3OsiM5LadVXa6FQjsPPWXX+/KR/UTbqtvTPqjJZPhnhYdrpD/nfyKob00tf0EJ1h8Npo/CrTQy
BgOfILX0kM0V7byesbbfV6rQzvQM38BWkWgVjE6OWXAw4Zb71t0OFMGHJitZR42nqmEUYezlguvR
m9lerI+G/GDMxKXkHiRRFgd0s8Dhpvr72/ADioz4GAGQxQycNAwDplNGRKa6qE5SUM8B2S7CYeQX
tEoxW485Yv9HbScvdTENZt3bxB0MzATMuAWhMx7LT7dutf4gvRgF94kQZqqC99T2Vq5H+/8YvIiW
R4t9SXB3FEDjNwsOEgeT4C6pMaLSOruXVUVn4LWzgaJH8V4MzE5USN0HIjpRTLODSdJ1bTEWI9lt
IsvRXoSo22SlAkBYB1/CaE5Jm1oBDwnUAq9VY6I8pm6RLDitLKxljKteLEiOF3eR9TLWEsDzKjLv
gkUPUJBCy8OcXmKKs3+yrBxqLKG/DY4bHVB/Ytdu6sd7WdVL/KME2kApqPoZumMYLkBQj59ESsKk
UhPshW4l73ItxYSaZnLGMBCqbQgB9sot0VxxXFtHI+yzAkID/oSuDWrBBpLWzZkXJndEDEwLaogR
ahValJIcvkCutA6pR3GE+SigrS0jXugbSwXJjQ0P4lbSF0bsb3SagdB6I34RmpuOhxL2LyaLm2sv
vjToDMGIKONVO7DBgp1DAkn9sJzIEKfLg8JEE06I74FIec/nfJQ4DN850gzC6GWp6X+WJqvkXMp8
g1Kru6nuepHOq3yVxeygPFfbrufYPkK6+Qemt75oLborkN0jvYqPjkpe8y5QrV7j0YzPJrOM7Lyl
rEKvPH52p80EqdxcpbG1HkBAkHd1z22Q6wXNsgDhz4M3BnrUa3XdDRV7BK3Jb/RcwWaAYD5wllam
scKdvK8PInTZv808EI47sjACTntpJ/u0f42eio9uJ++xYb2GsU9ppNj06EKZ4mKcZg1MONDIS3I0
FucLItOy1vRg4yuKbOs4W0BMrIZVQY7B90lLBigj2tdMtg4EifR0ILAZ+RV/aklAre5gw5nbPFXI
JmxgOuwhpc1Cg/DA3FkbSH6rUu+Yxjpj2xq0qdzSYMkt09mEANRT7L9sXXaZB9DB701XaTlm86Pc
12LtOXYw6ixQ27Z/C+YWMyQ3NUNrAHsvh6jICwxmAb4B1V8FiZqq3ZzV+wA/H6pw8fnMKBS8EhSB
yqgLGDnrrxEflRUUQknSYkXkrG7yySCaF4SHJujPsnx63mKALb6aYI20UrDB+MlMNla8+FS7npHF
OxF454GfyOjd3PSxIWRl74n0byXHEzXTOar7k9nNAZ4xT8b7DDtAguEhaKYctrOIcsUaZwNHSQhu
Rei9dnk/CrO8qTIbwf+ADD0B6B1s6ArbrEL9IXU/HbkG6wekWI4llRoof670dZ/9lyCvvVzevP/X
/oJZqttaHJlweelG/kKyJbCRZX4y+M3Cvn1UdEphXEYttiUWk92JC0A1asK3sXrpJVauAJc2OYVf
OI+neV9n9gEjfWAw/7I9GM1ZNVDP+Jow9KgNnBPBDoqL9Oa4PgwZjyD1wp0vepQvh3FETZ6ZrBLA
lXGokoHhG+E4/8wzwiwM1/8mtoeDe2ui4ucnNo9AAYkM/vbUMuWwprNkq+FNOnsz7qsNx1Qasnd9
GIjC6ActJZLRTnHtFmUYasbgDGxLc3KLcpCTg6OSX3fF5/oXfBh5S5EQ79Rc3MXE8wjG20FYGKbn
QSkJaTHM+9uodtQ4/mQQNXxr1Nw6C1ZkhM97299Te2R01xNaTJ5sr73zY575WGlgWMRDlyhBDIIc
lka/GoGkNWKG60dXg9Er6ILkNY6VP3yQHqVo/FaILleLkga1StVMocN1XSTetad9y5MZeLrtV2p4
1yB4ltl95kSHvYVmnaeEoJXSvFX/INmsTmtZPszEaDyJeYruh0vBdmzOYv0EXhmXDE8WFUYNvFk/
BS79wb8zQkKMWMY1OZxi3H//rz/zrf5tIMJhXa9sn5H+4ms9FVO7if+TIO/1soNphB72D71YnnLF
MERKWH/lJq9WYcfsCdbFn5SVrfPgvA+EM0gwoV+D2MP72Q9JvMFryElx0KP1DyhbSLVC/geuqkpc
s5SlgSnpDVj/0oau5Lr1SoOp+mdp+UTyR6i+U5mJlguYFh6UljIgR+kKYpUb6DXD/Fh/l04dW6it
6Zn52Or36uL4LYRZZba7bqtN210R6j1le43EcDzUjNEGzct08FgPb38Y3YdST3SI5mBVGzSfqp7Y
E25j6+F0ICpyx4BDnmEtLdDD4g2sF609gdvrVFru8VUtQbt5gdezkQqNFJ+1NlWse2SolAeJymSv
3bvJX6HDJ664DZMAfwskjC8KSD/dPwwn6GPhhazPsKFJc5vJun4LXH165NMH3NEoSob4IO7peqBe
0EV4P/PxyG9Lx/exTsioee0ZrJSLvu8vmudJZbrqX9OeOSZs7I/imcGba4SxR60u35fLdig7p1A2
SrdunzKSQIdDEd55maRHbiWOOcokUgDV6j0sAf5QwxaqNH0PsmuKaGo9gY4MGG/zv48hKKJz8fsM
YTDo6c5xPVNKZ2jVPlpygLTfFluNupsNpVj3QVminOpAGia/BeEdt2qWU5hN4ZY0iwjNLUvn9m18
ybuzOwDyC1f57axDPrTXAxwjMbuhnJf1P6WvlaQ/z8yw2rSaXR5EBV8TCIRZKY8LqEutdgkX1Klq
s0N6OHO8KZFfXN/KuCM57yqJ+YTFWDPwnmEuJIqXzEH7UHOYGNEx1lr9qS4BDpDgWFOKR5j7Id+X
Con9oQgOq06co/BbsiR23TQCxr+d0fNzWjHIewK9xsDX/PvPvS6MGEC5w39qKA1cyz2PL8fN/0/x
U2MvQC30ZBLbNIP2a0QPQsUvBKEvxPLP+fs3e2yd7n24EkxGM/KUe7N1V0RUthPKlgc9QQsnw12A
FQ3Ra/N0Jz+g93V/yqZzAq9zIIbFUv5BSAQbRpAmlzR0EZAr34qbn5mvFb1jqdPaIhHLHUgVr+dh
SGDXOs9D0FHwFaFp7RoDUYOPNFkRkz2MC4qw+04RYx8br2/cVPmtoMRiiYyJZj5Wi99Z0bitW2Fy
d3Cvkmq8+hxWNQC47teXr25tzNLRYIrEfVQZf+jGmvex3eFrhOTCGIdKWSwwhx+sRaNa84Fu/4kY
jNTe7BP8F3N3mqMZtBtY9d32/elJXDpyyUSzwBkOlB/zkkPuxwAIaM0/oQuWpNTI7DEDubvpipuK
tRl7OQS/FRVmFyssVLuIgtpzE/moktE1oUPB6ubqod4hQTGGPku0iV1YZXPNz4rlLKjF8WPoBAgL
Fc6tL962NyitCd/zM7kMcpsFIE9NJb3XtvPqZbO6WpVNqK2b6RoFgjS3O5dQUKJlDmyCVKRWwJ7n
2mi9g8406qqVbkeGCHsyMjEy8xlsKwbCCTar5fmMFEdq2fTX6ro3nxP8BjhuBRpr/yLEyKJAC9Q+
rkjOum/fuq5/SGZC3fjZ0F/JGxKcGWptLg+r/GYFA6UesafiSrRUASvKUxEai5HNyTsj1UeDj9mt
eXKinaCWtzMYmJDNSumXQoiNFpppv5VUfz1EacrPFZ5m7T3CStu0Vyx5+w5N5d7UM9irgniPk+uw
LqNtwWvB07xoWJ/xowrlPWUsmpst6hep2TYMMvNYeJZJ8Nwr/PnoBKo4O+6HVraFqsJIvWoDUXtU
AIZ8dTS3Qa6VmPp0rLAEScTQPlh5osPzikRWk/eprTjiNl9clFtIsGCRPyJJVN/VMUQqd0wkN6fJ
7UadxoRP6/Tnkj/x6htvaIDIJ5oVT7BmvSGQM8nZzXt2lmW6lAGUCyr5Ef0TwbuWrhrz+GS/0Tvn
ODfx7WaXMNuTWVsH/5JZ7EQXt10QV80Z3Ea3oT0SHdQgEj6nywuoumWxVDRzfO2czqZpcmj1w5ld
lFuz2H6Lma5B+F6jzOvbVJLGabCtc9cu31a5P4fQi4AHwTbE8ahSDR9NqXY+lYR3dLteQVpG8IsL
9VRyKIEKtuDqbvcdK8JnTqCsEfaS8fjndKVPFW76FtmgffDPWuNp0yw4hrGDNCYv7kWNvY4OaWSk
KprpcQM5pNneGqD3EUJhel2M7nPK5aJGHpZK/QPzx10lZE7k0ce3nWcyVmmeUbwAOAH37Y8SKpoO
VLVfs4roNYwIr+qV2scial4wa/8NA57Ux2a+ORoNrpIIDIiRsTr+cuQtsq2EPfrj77o6DnbvRzZI
Ru/ro2MBvnsNejRW0vOCN+TMct9QCdS02v5ivEyTY0NzyZ/RtALNviVabruXxUZmPEY8RHztJS1+
xZ6KD9VDTKiirOJhJTkIcPxu58h45Q4hN8MVZ+0eLrQNbVIri+Ne0NejSH+zSSTev3yFegLwMcJA
It9jDowq5OfUT3EIh6qX33XHPqftVMSZX6mu5kkbPdtaPffRY+ZjG+8CIwXExoirFf8qfUtRKqYD
qhR848jg1YMLQ+JRF8x/UkpywpfCh8HWOzRqgscck+CwHhGcbNBhvK2SiU92PIjX4hD0T9lYfc6M
WMs9xwjwoIJqaSScOSk1OLD4IGmSvb0uCimhLd4EQplu4Jxs044NQWYf5b9+EHLAr2y1JZZE7y6t
vjMDwZu5Phs+7m4if2pGrvr9pA9mTB+qqYnxkhDovw152aoAF3JkgwSyDgiJUv6a/gIT6dQPDYuG
R9B16RaqFRxNKz7M4jeTb+KPmxCtESExdYYx+BiNHDL8PrwQ3wTy5urfq8u301mMu/GmV+QKAjwm
ssfZCJctSsZSie0O8i7IAAco0QKJnG95cZ/UmUsTo4nPexvf2kTdzHiLd8n9+YBhCWnC72NvOBjP
wiMghCvmbCTH/kI43nXl9EstMK73EeStRStRJpEJFvFQib+sj4Bs1vHYMjCTkzFsrtoPp6cTVK5G
w/5H1WKN1vfLWV98ZWYrAyMwezfdXEjJZbb71VNrjG0wZBrC0iGRT/TSLEX56CKJG1G61EDV59cJ
zwVP6wNuP6R2xuDx0jyR06U9dWmVE6IpTcz06ojrjI9yj7oe9XlCBjF+vVV89eu5ON6qSeVoy+FB
VrtDHxGeOUa61AMvfQGt+ctNtG6OK9SQTWFhLbkHUBPQI82PEzADvDmD951+jnngclJLqeNM5wa+
V+3oa9FLssIR7AD7C/9zS1D56z7SxBMqtqSMLMAxkEIHtDac9cZXUU4McFrgpeoW9lQK89+I+yXu
Lp4QJ0xz1TeNfrsETSnSlIZheWz7Va/nb1ysFwJEvzPuH9j0RkPzDV5h3ZvyWeWGla2y/Nhp9ZvZ
f2KtitpCpQLgrxopWcHn86iDULOfgJ23RJx7nRt7pV6p6ALpgm/fz1/huzivexpTF19tVKo5df3V
2IfYcBv8T0ntoQX6GB16g1DGAOhooc0LBVoKZ4IklgZsbCACFY5b2dshJtr4qGptMo4NVvCooUR3
GfyoxYNFPMi3tj67Q/+krSz5TPOh0przD2OV0SaSCaIy1WrwytqNHtXgcys8BiLXRpBI6jrtjCx+
O61vFzhz6DH3bPrrVyd2pbtEUjpEMGbOeZANQDW07Haa2+8G8F3gHfuqkJgj491lFwGWnZeVrQNX
GlwgV3bLjkgW8oF5xtbpODvG8GN6A2O8tj1BzsY6HhVhZv/374nYTClMWybbpuUlbtiEQ4zG7EGK
H7DcrQZBvKJ1mnrHZm/bxYCRbcueOAXQe2BZrYELwOXSFsy12DkpY9ouCc9QWpHI1ku5Bc+XQFtM
S+zYbmVAn125EeGYa7fbrIAV67AJPS+5ygHvaJvU3gOOuFL1O4rhg2J8tjk9Aq3eHnVoQoQghqVf
XHK2tOg9PuywXvOJWTuWVCH2ZNKfXDxkNMtZL81l+APmSNPT2e38PnjHXi4ppn2t0bxIt53aUMVh
beMy+yHDA9o05okHN2pnv+hNQJmgu9aPCFn2PIVyA7SLGP64iGCMH7XwanJyS/8lpQcS8SyPxG6+
m65L3bxnzG6Nl2pKmOYnNcu0rFSsjQg6mxvrM5JSTccDTSewB5CZDvit4+PcxC/vDXS6cDOwSYf/
U6ojMaBMi7iWCmgDCUaGsfdeJffdqMx6gLLoEi1dBBe4WNQ8APr/gGQJk2ylUtJBBK9Q76XxCWun
UWKHDLeX6+Kv2OiQRPAKYJ18VtwRPiqJFAFrP8vnDffwSLegkqibXn8HNazDV4DTibuYckHLz+wQ
aR0LAhq/j1Zq3/McHuXbwktbm/xoX2ox+qVz5i8jjqMHzziDt6ON9CTooKadm9m6T4q5nQH65Xd8
7bDEVPa5fbd8z1p6gTy+9VKKfSmgKQ9TWgou/jv1kM0WaXRCWaIcpWzJVAvZn2ADaOuE+mnmXV/P
5E9yCP4QMp6b6fD3UECVNSrtsUP6AM/h/tg7giqng87Q8UpNaT0Rd0rcr95HEdjNQppS6Vi4y6bh
a114ccBTtM886P2ayfR/U6jVDbG3JWHInKz0byvijaJtRBN1EjfsXt3CUzubf2mS35MmEg4UeZm6
ZqEdHxAWOr/Gi/b3thFHIkPljaffclhUWZkgM5IgMvq+K9Tch9EQ2hA56adIWjiJTtuXdGoO6BFH
L+aWsyRJenzNG21SMCd/7PWIweNUZ5q9BCEgv8klLz6D2JAKKIkvmpQ8yrJWBW3xXxF60AU0tUR1
WTDkugYmHCvGQT65GC8w9UuHEugE6XC71vpmtsQl76EeAkT2gnqRkPOc/R4DqCmKd+27cEo8Uf6l
2Y3zgcqUOXEqYdg+L8Re/wM5kFNJLb0iS2WfV0rkcX7sgUylswa4Ea8tLTklZIYGUd8ExiRctS1X
aAcC4aUkyQDszFFSZlCs+y1e+1t6lhtOSUqDJMHLgqUdYUV9ERH4rQYvzfFgYKWnh3dpXqlp4hrv
WoszmvmUi/nV2T+6K3sYOoXgV9W3KT29oMnXCE6tagXXN+nx7puuyETw/sriqQLaGx4Qkoron3qo
/RXrflJgvRl8FwGLx2V7QdsQz9gXA7VzvdcLEK3gj/sY/xV/80YnPEciZmB7SiRsxPPUo048b818
84sZraCbvD+Wjb55mgyqeDKVwBu+CNWYLCFWuV3LV0HXm0VnMJQA6TV3rmFLTDZ1ZO7oA1w8hAb0
ssuYI+q5fd1CiO6nC04BIr316C39UtE0EX6Du8Nc4xjP1rzY88SNAiDL4/7GixPhvEphlQMiTCPH
so+E2GY7jW1sJX5hMakYmDPmUnccbe8PS1dcFugpysJ9gPGqWTcMurIRPrv3y63AdP5pJh+Qw6AF
HYIwJVGZmuTJayvWZfPo9YXeShNyAu1qyPKQBrKk5xJWQOhHduhRfHsWms8JNtAOTYz+xGFAbZWa
IL0WPGdh113IAp0kh1zmmrpQ76r9hGJYrZvDGRLdCxoorjsllFUh7H3+XZ1kHtikzFl08mgk9gkm
YnS/ClDGd0h23s/MPHdey75oBuWrpvJOiP+Cye0AcWv0t814DccrjAr3QtyPQxrQga+6+EsrjTZ8
3QSERUbTZyF8W2OS+S2zPjyCpyVot8X4lcPJk/y5qJJ0zYchkhFKZXjKdOwSYlNs4yuHMTsEYFy2
bb8q8RaLJbszDlfP4dGbECckRYX6ewtJiiJQ0iswrvlCuR7KPeT39nb5OZfFSLDsR3Ix7/8nyCjD
3SG5LBWb1LWPLlTNhdD7lAZCQcGfkB21nmBp8olm1QzsF2NLju2YjS/nArqjGdpXowaS/ffrqPuC
PamcPCLXEMWyOjqc+j/5uxb3ncXzpx3bxjgoq/nGf1qzZTET+cPDsyjVpnhdvfj7/TMVtAgYQ/Sp
dHLHghbkHDEeXkPI/xvw6u0qP4wbuz6dCLaAvoPssMEarI9UKM0WoXX7iSvfwSQOYFRx5m0TGHeJ
0lnEasjha8A2xTOcHlGnyJaqJfvwEd/Z4ve5MWVI49gryM3ML+PlVfsQVWWS16uWAWJSTi5V3hUj
s0gbuOtld3dzXI6M1K2wwS2+kXi3jflyVduAEiFXWPPQidYzPFjZ0TN8d/txNf+elWYvoVxRFbNe
LPKnU7jrQHPidhUvg2oX6S5mkuXZUQmib8aOOSkTEEM9TqmvTgm7ODL0IYdrpyUg6jwrkcz7wVqA
4J0ZMbl3EYalUhI1Lh556nIV6CacVCow+glqUUZCJqIci1KGmfQ3TRNzNxRMJkiQYZJuI2b3EU0j
KJONHp6khWee46y2nLj1E8DMWgQTCn8IU4KUUkYZCqNVoBnsb5+lK7h6BfPyUtbOxKdXIbG2IxvC
kgx62GTaOPQ14upNCBmt7l0RMHUm4eoyNVVEHScQVgZYC+bk7bCJ2oAdUPIcFIOVibba4mlqafAu
/wDTUhsrN5cAuI0ooMW6r5KuE4ZtFkklMk1NSDRioH9L0yiVPPtL9/akzYKAD1w0h3L34d2ppBow
hcEFWKsyoGr6bt55JrrGrxrp76ueBHqFTActRzeV60MzcIFXyRjrpxy4PTO/J4OlrcHx6dky/ehG
4Mhc9p81rX4YOF8wj72qWFgQG1v77+iFiyN9Mq5KtxjLx373euvUMAjtmuYQWcyxTnxA4Bg/APUn
pT/CsE6N+vhucIhjydb1/JYlDrjRoAMXQqNkaBh5EDGJy0kR9JZ+TVSiaEI0c/0PI3MgPdJ1fC8u
ojLbQp30vAKbDYoCD1wOLuuM8HpF22MeXeepWU03MgPM1TP3G1ExiPuigV5chNnQEAssOTe5jnSg
V/WbrX+i/AqSPZP2VZLjIydEMYLJnB/Wi+grbI2I8+AqOzKS8VaIN95FbwJ+1L6KWjzG+bDcv5SP
a/co9LetkJYlTBiFJEO69Nm6SVgBtTUOtMvIjO6nYIkrwdLuHcxCjFnzqDlQCo16DQ+Xes/BHQTs
5qgtHYQYYSW38vT66dM4zqLgMrn+vgARsqDA/pvwDGt8bz3sbVSMCYNqNZU/2Uy4hbFO8rYKg/s3
munNdeYSovp9g9nFbBplbfw/Z8ydrL/nBOiQmP9BqL4YllkRBRJWjmcYjNchJtlXBDhZFagmjTpv
l344xo8jm+g9Jodlwpi0RPatZfPaK3T5N7HivaN98ava3GEbvos2Qdv7Ku+Kc+/Vg58rvWwAE+Ob
SUCqsFk6UU/jGN82AGv+wCjRxZoqI0ivDHDXMIDC9v3BZPH9fWTKXfhNjFMQpy4fVL7Cun2GVZkW
ZDVMwoaA/yIP+J0WWwHjvOSR/+so2k+C1ygwiPvtwL3gwIqB52MKId7HeQfl5DLYnehGxxv0PQ9p
PG+9xIyld4LRVUzfUngvJm16OZSN0bBkmG7uqjLppXPNlYDY1bCe8HOKBe0F7kNq37lzsf1g3JvC
4kmWKU1hva5pz+uqqprgfn5q/v47YTXjWF4LL7lOOB5hDmh12GDPgOSnw4SRPHxKdaDF1z/h3Rh4
2RpVVg0T0k/72FrJIdn3pu6H9mnt/776U+hKY6USML4EFy2UvRSKIxH9V2OXvFEksklsxyzNdof4
uJPuJfsEBkpU9sJOUZM8rOfG4L6TQyCFVRIpMZzC+nnO6rsYSaZMpAn7K614bVQPvp0LMXV0tqCc
ONY8ubcq41Mv36S5TCkOUDr7qud5OMjdZbww6t1fz9lgQpcxZoJd1NnNLxBR+NucoNfgnLWWzIQe
UYetlO7c1oXF4yREss10xlQs6B8Hy1mvj00ZoD6gdNp7xojDClU86YjXyH4ggHBJ0u0ubq9kuDmA
wAdCJxAve9QVTSL213RFw/dQzDuyECCX54mvjM3c4PGQ9INTps6+THLlNMCvwI7EYtF/Z8Qnl0rG
N3kBDAL/LUWKy6ss5TypZBC/mOi4/Tegh2PLErvMTyuLgTQB38gVnjxVeUMcy2yt6LcbpNJIgf4u
VZjSN30hCB9JRzF3jlay2CCJnPctkgXZgo/QBmHDaZLeknJl9KDwhl2Em5MmV5aiIQE89ALDC5fK
BkWRpGjegQdz2m/S7lQZR8zOWN0fS4gEf/ENg9v2k8vQ+Uq2KrQsg8JrMEz4HWtD5uHoVs2MSgn7
R/JZj4dzGPtK+WXjska4pQTh8v+9Qf1FLNlPLl1V2wzNZbIQ/vHL5G5lavq5KosVcsDgFK62AxHS
BZOq6lg2Pxu0UwrrcsChIwr1FBZbdlWkmtgKYDPulNrUopHGKVrUUBjwLwf3+TZV1gG/jZB+XCsm
0czqkWBFbojgL5kGo0uWpmKE/PlkZuniSHBssCantGw4p6Hpu08A8JIFe9HDZlsAMmMBkqAwfPzw
VUOCGok7zZBmTrZAFFXILkwHUBHXAYd7ejFp/SFINd2Y2aIu9TYauFP7PLNXH1JQuIfx3mUAcpNb
N9ojmfHCgtGg9Sgc6pjIYwQvcRzcExcIRtqs/DeXjaaqLaZ8q+M3Sf65vEjrJQMPuju2vkuFT6Se
a5OlWFqeEcu4lIa+RhiSQYJIN3i5qdhFIf3kQHnIuFa7+tnFP7ndOXrZoIAD6NaoDMT9qOH326Ie
KmmHjUjznpRzh2sh1zcTCfE++YOvqdI979OF0NKtdcweXv5VkfuEXtOwt3An+HjOjqvW/egWKuyF
MQxq2Jr2Z0UQOltVYgrTAbTsvQySRN/eOJ2Ipwe4EMVgboxwoIDkUkX2rw5qdZAnbKHhw3ET2EiY
yyZVMnMv56QfkZJJklKR2MDswm4znubZkwYjjNYBP6RiartdeIfANTW2GL1+vIF+XA8Nbeus5hCY
jpJFdUEXOnI5PE1bNSbt6aPp+PYUruhWWJiVoIEEhX9w630S1A5+h7BFkx5pVPDAYBODs6w3JQdL
5tzoQvkcwtt1GUscOxHAoymTjqseG7G3pe4m9Y2d/dLdykevfNh3uP68leYWOSBp/5Eo3uhPek/8
23paDDe03jwLG+OC22PU4bsDGMYhv133GMaPMhP522fxbVJiMn199ewqqXdyMbMK3hiDe4i0tAwr
im4GHkkiMkm72LLP40MmhvJBTFDQUNLDWlD7KkLGsD/HDBy5nw8+n2mTSOGqNaWFkOS/esELc+CQ
KUx8KeE4QYO4LNkSdV+N0pW319czShooR1FfsOxdrn14EtDkkjhO1MwE0hX4UnzBtJFKp/bcnVkP
4uANb+IwNPgRxlh8H8PLNPee4t2djc5y9gT1zLzcR2xOyiTSX1Lv/U/6ao0L5fO4tLnXnXf1SHP2
31PhCf3k9J5vYQ2Piv0v/KZsltmmnTZTp735VnCnaLgXNdJhKzgq9WVLY/VJpPWXY7SHQz4VKW7/
8zH98kj7KPk0aA6gEDWoGYZb1um05Z9cuUopCaRDt5fkQ/4r2qWUmMSljXOU0ilj9e1KLg9gsjCH
G4a78ymJd7a96oG8HmN+WXG6r2xmXauBY14MnUnabY3+z/8sS0T2aUh8G0gWRviKX+Ac55wWAKAZ
ZlnLCrwQSmTcJV+dKau3UGdbfj13y6S6JQw+wmPzbfdEPYBXcRPABCCmXATWSCIF6czGqNW2Xfiy
yWNraYFWaZiR8vgFJkLkyQQl65WyE5+irNWXxe3aIABqFmqqdUMbxxf/CjZ3HKf00wJGwmmhk/aR
lf614rG4DWdLcXg/r8Uw9KorNEEkbnYgDPFMCMWNGYwIuSG1m7ZNv6diGTSJ7+TbnmIh2L7fNrGk
KfqJXnW2BkNxE4a+qq5xc5p5+Jb95k7d3V2Lc1/wO0t/z6/g8iOP+rfNLeBtDK7H4T/FIrsHLdO7
ijxCBLuEu/uC9cnnTcxaJiGzL5Bl7F6nuqU+qYaNQ9zqpldilQqIYnavvtyjlzEwEQK8DVpMh3OL
yVsxf1ESS0IqV4hkismn+QIYg35teyrjKfp8ZVbVXENWiVyFYbzZoJ0yqfZcaFdEMqMz5BVGyLgh
QPuaz5adOg71mkJj9ue2zmlprMhfiN1Xf9xmhtAwP5wPt4UiFIzQ5zPbrXfF/2vFfwhCvPQLvNa/
Gjb1zTO1IaZy4zxEdFT6EZ0B5Qj3ChM8Xqk9xmDWb7KBkumVRR0ejRbZTvvRWS8Fa2crFHhYZ41k
rM/IgvgPXBsWnPK1bu04LoguPR6GtRwG1o1Ob5dGZkLg/39Wa1TnsTb+qFJAxPP9xoa3K2dmfo4u
q7/aZ2/Ko+u+s/yr5wdGXdEx06MfAZUoETNa/Oq2hOIGowlVFnAluipJPs3n0GMhh7VTminwNPP5
dYOE7H10A4bLBxEgo/AWYc4ADWpRPsJ2UAKwh5OkbD8KuOFGwRZPE4C07CNTydAYR3rHpALHj15t
1mHL66mADORloOUwib9kLVwtIOunjC1MbUmAptG/uibi1GNZaX2RGTWwo8iTnkdGL5ZfADiMkuML
Dwx78HtzzU/EWKC2P0DGrH6TFv8d9qvfBEAwuNDig36mtgNRH6jd0ieVdLW3OMgvXe6IPwOYXzLw
wX3Bxj6xYQKpzCNnZ7nvmBdIh7ZqJ6mxgBT09OqZZdgQ6tL7S8lVqIFi7/y3I7T/EAG9KzjeWb2k
+IGT1QctTXJAfZydDJ+yo0xpkyGg/fAPCH4SAlYaWwTS2/Q95ULsJZJNWSFFHB4pxt2xtRPQSPxb
iWbtiJpX0Emx0VyclaLNO2BQyefqsvwp1iJYGRgiSChplZ6MmO6o3plxZ1tgXJFFiD5S9oG8JQ2w
tFdcjo5UsmA//nrbqlfzmZUzIxRWktOwgMDLYaHx/GzhbndRaPVP4Czxv4xODpc14IGnU+rgGwP+
EFUL5MfavnE9vuEhcpQFrzGCAAOI2kClrmeqTEtug+QYlJbGbuVrqujS1xvL5tJYTlcVOp0w2CY/
HjsqaWeK/XlVHG0FPD7LxC0b73jkpXKOSz2XGqw4LbLMFfsDNtvbxa3dWg7fFJdCe55Xwg+UJUAZ
Hk4J6mq174TBA+wNFvn5GAEFwb31s2kraTfwxhssdlZXB198bT1ZOAkOZV4tTIswtu74Lu3xI6bN
x4JvQhFDCmiUsyc6ve7cXSik8DHKMZ+Efou4BtMsPOfs+qygXk3jlPKv3UzCt4QV3B4YlrWVqIl/
M9Sq0JrIXEdGgSn3wOK2GsJiUVKbB5W/XrKz5LHom0h8gxV4hpPKLR03Ox0rzpukpnz2lJV5bopm
FIrnNTxl44/vk09vnXYeen3GQ7HV1deTmUNgRaa5HuAvZjbT8lDYre3bDwo8YJztNnimKId77nQI
k5ytugEjUC7uyJqM6q9StFPjaPaKcSBjiJ1FF7O6GIfRvMA0uOpukUycVzfjmhLk+ziUPTEOMwCH
Zk6FmF/0I8ew8lCHGg6y6FLqc2s+/qaqnj+ivXXr6PUVEEUhsE3DnXGWKUGtDfFu4Ndvx0a/c1og
SpGa3n1K/t1G/T57X7P0JgFcqOItAtS7oaH6a2V5YOnaMOvGZfyJOf1ola1nw47RdPDmDfK40Oan
Nqi3hh98AXgUKmyfmof645ts4GjeOjfwiNJcrJBJdNPKr1s4g8CVGNwmP3BgwM3xmWVKBi07FduJ
JRCyjAE9R5djk2rfbHJu/MPYaFs7JwSC9KFXacLjE6N8upTpth8gNm91m6nsp5uX29REdQXivh1j
Izpv7bsHmKWMeYuWhMlIzoBbRkM+y7RmrSvWIhjyjV8bZgzA9AMtmG1nnZFofjCHiAgVZCsVI6N1
SXsbylFsqnOfQu4NJ6tyfjDFRbeBG031A8nu2AlD2EwgsHd2SCf2BwAGt4kSA10ZND9o/f0S4Hj5
LOjx3NmgytOclWVTG3/SotnDd3ARqJOQ2lbynY+UZNGluuyOG49WCD6rVg3M8qKLCqbhSa2NUoko
J50L7Ro4Q5BS8W35sxEF56X7QoSYByv2JppqR0qeAWvHipQG3+NIu9Vvu10S61V0Uy9G5Z735Q7y
OufiPoChJjQGUACEJXOMe8Z6wKB8aggMuStWGmF5GPexI7r2M+8rMd4hN50NA6Ee519svHddqhmU
ONYkPr/WDyl6zADoTI4I0zcO2+4sO+2yTFHRo0iTjRTs0q4hLXWPxc5qxpqFgEGJdzyLYRl/yyNQ
Ffl6Sp27Yr/ZrRbu2luqn4WKc+olJxzfTKderONhlRxF4sD+FrYHck1qCDDuzwfAX45NDxkBmavo
920ukTytStdssQc94aJzZ9Q4k02SO2ItCdxA21mvvJDpufciOsk9qFfDhj7XUQ8TJAtl7UXK91Vw
ahZ+JVQv2yELWUWOznSpUyGENz5H5OM83sjfKhAATacjnzl6EX/IOacpiS69G5hv+EhAbgxr40He
Z8hGMhMYcZk9lhzgVW9KBEZhQ2VBVHbi1zR2iBvzyMmBqGoLhuFpErehQcO5TSWf2ViQzTSxIbfS
FMbDi+JXMiA7rKeI17Acv2dkOzFe0daNpDTs1AOXSNKUFxzv2U/KJRERROnZc3WenvCXxockgn12
ulf17NyZMBR/j0z9dd+1wVPir5W/XSP1y/AiCi+YxlRc0/Mo4Oq1KtNrEMc5hSglyJp2YKlRq2CU
1NB5vNqehMv5oqayB5fehX0ZzlXFSKaJoju5Q+VYaGkOyBYzL96qmaiQLK4tnccPdmCdqFk6Aybv
H5g0b89zp/MxLvfsvrcQq9f3/YoRjmdCwPzvZqI2AyVoJWFRK2JDloC4DQlqzmLM5OWHfbUKlinZ
OkDWB7WN2nA0bbu2wgrGTqwvIY7HkCj9Y73kj9Y5WwsT2b/8iD9CmN/alWpDtrTxbNVHO5P6Pwz0
WBRAlsNlEcTZYlOTFMYfWp+lMXTjELx5KAB/1+zrs9zTQCE3pcxjl5KFmtQ2SjHZLSA4Rlb6DjPX
WuYKGvyyGmWLj1jeqr51WD/YqmxcX8E3jJ6JXaXB10v1QMjBFRpTbkb4gWKQN1zwl/frjxTJVoUK
gRZbV+BSfVPA/hfQWpZH212X0oxVX7cfCL1EMAKfgtGNzEPdHDbCbYhg2Sj7DFAZ1a+wxbNYOvyj
F9P6Kv2k9Lq4dTh1zRQwHHwDnARFa+ZoQ1riNrRbmKtRT6WWM+3gyjMm6OAfTdcydma6KCnSbVKS
/e+B+g6oyhewiGxbbmbWSM3k/4NMX8WXQTVypnpYHHSF3Ad3kh7efU3eFT2NLNUhZEePQQuabvlG
YDoPYNjqwzV6R4AzFKj7Cv3JkhCLatwFyxeQwV1dNhc5gKS1CTlWxO+NlbQgTKk8jLJpfnX7ylxJ
9KZlGwYef/HvatCn9TIbDzErujzNc3QUF1+vme5tKtYMbNCwf0f6eer9SwUS/ly4Q18jqK1U3CDB
AYcymztd+8VahYqL+okZO2JAR6LD05It98XL6qNi8jgMcWcpb+t92n+U38w0UYqSQqOttzFfx5Cs
OyVTpomvT54Do7+kaWuj7U91kNgBoxCiO1rrKf9zG9Zq1wkyiCSktNdGR3amHlmzC+v/VI2MjRK2
esMoI3Plk7NDAoyuNcOhTCL8g1eze+5B//bp8rmCheEEsitFk6b6JLsncgT+MltCr5XCzfEZykIS
LvMMk6LYVna1Nm03vcuIuJ2hgDU7RN0doNZ9oSNMekiZ8tvHXtQnjrHWO6J4wsNuQL2IMejC9w4k
EIGN9G1bVh5MSd6XU7Z8yy487xFpCVqLOo36CEJSlCwQRyGLwJ5GkWjsbfet+9LvDPD0Q4A1qLTW
RasEeuFJkSBIbCoI8IK09Jz+jtQZbx8Fj2eV2Y84srKg2jXOh8+4/z6XCTY1A6FIzoBWwafth7qT
QoG/j6kBapNh2UUFRdQdELNcOw0LVQU5slRVNynLx60YNGCChltt6/XIPx1vreZLVWTv3+6tOrha
g7cY32CUjr9YhLXUFooZwvzrFDRx8oK4dmijxjAy5p/ZgTcnhjxgQFUdLUfOBh2cv6LNb/2/STYy
9z7jpHtC+EX3UB9z9vgykYSSw6Xxa3Q2k7y6z40vBpHmaj0Gqj7npu5K7DNywGAj+LXZOFt+hJ7Z
bPEHV7FR0xDTDYXLyFAp46jDLdLUZlLMk/2bC0Cp50NFYt4KXB9zhS1c8Z5Xwn3ZX1MiKOzFPzsY
XH7h57G2ho8fnE+5ozbOcrAqyNkkc6BbHwEDQS0r4QsN2BZECzSd9ikW8px5Eo6L3YeB2f/OCH+M
q+BPGA/hkZhsXdsPD1wfYl1vf8f2KzFJtN7FJbMcXrYxYnOghdCrloSkRj2lUjaO9W2IXYW48ooy
zwAdJAjmdy4czkTwPaIC/r9qIPPE3uyHCPA2S0VgK8DpYbxsHwO35rFrC58tPphW+CCyaxicGyCp
QmgTiDfzx1zdD4nPTBVWwahyXsD6iDPWBkuVvLG/66MvRhovpitmMZRlgDI6BuKHfZM6+Bnk6xGV
UNSikFzUs/Jx9UUo9qSPmx1jOWjZFkQfxgMnRsQpQPBURGrMOqqNlZ2WY6L5obnNfxtvPClji7R3
oFEEP5uz2OfMdctW/+xl+7Iat5zhjmAqLy0FxCTOyNV9GnBpEyI5AUtUcsxiimwCSKTFuXnDkl/E
Qrc5VEBDtdmvLGj8vDII2Pdy+3vaNUPeIvvk1sbCy7sB1rp0lSHNx8WSAk+ksdeVitiKyVizhPRU
PVcFA+6WBFKkLKkco2h0VglM48oZHurENpCFVOMrXo9S+CS2CDfQqevSMDs2gA4WmwojfxEy7I57
0aYtDRkID+KplU7BT5jyzteLU/bwQcJZoJ/kxFyX9w1Sxc+fWH9N1R1CjYjRSe5orySr9YJ8Yejd
F4oSJmVDI64FvrO+qDh1iA5GCaUmcQm5pguQgaqYBC+8Sz2abHcMOvQrB5ashaFK671XN4stbAjQ
bb8pFWbKD8hGuxbdO0tGeLZ2eNxv6w54gidN+9P+0kAVxc+SJt51BioTFw5jaN/r0CU66QDsCyf0
Oidm/7o40G/5+FnqehdkSzLb3i52H9eC7S+Hd9DU7bbF9SPlRdB/K/QCE9a3W61Liuf/PT6nw63S
TfKl7rVfg3D+Gmmu3CQ3trlFwPm4fVbstVW7iWQ0vYXkWWmXeoknmuMoOYPP6QkdW9YA1GVfdFxI
BbaGQhMgdth/dVuCOZ22Kb1uV72CnDNxZKS6PrYQlVwz/pgQXXHENLRtddIcWNYOkfHsK91RS5QA
IwE4Tc+b/KFvIEM72PY5oLThWSn6yXfNXHnFssDx5vNOecvqImLdDCDkscH6XxrXgqd1xdQrMbsH
2aXxM5iSkKmPkiZV6q6ihTo/X92cmmdQ3B5sR0Wh8cJnTMPO2KV4neDSkI6fcu4Jzvn+ePuP1MEi
WsFRlNqDYJhPUoQuodkKRlwq98arG78gXgEIW3PgK9PdJ8WwsKoWaeLI4P5raG7x5h9AhUzo0tec
Q5i+W9O9uvcVNMZzRHgF+CEb+7O1Oq+7Cw53DqVwjmrPGI0VjVzn+zGjBt0e5J9/w1B+LDQOve34
I/pps4h6wb0zdjRuQjZa4zC8AOKEIZvOjK7+WMSG1qTfw2A8/o3PHs6k+b+GtNMXacuJbF8GgrX0
TwZ7VNjQurqDpTh3jExOHw7G7otbWBbfjrXs45YR8EjF+mLEErxh/dnG46Onk8M5mOycphrhn2Wj
Y9MohKTUXAkKeRoB2j5aOo1cYucle8aONhgWTfFdwwj4EEloVTVv3LWoUmpkygwRyQbqVouVuaqS
Zoq5bgqzuC+FFcSxmjQ8NA5kKZY+aPKNd2WlFOsUnFKOtJv9mcWcwaBv9hFwOXq9UmndOjdevv+l
kVISejWvGOBZva3x1edPM3oYBn9pAV1pQD5kwNFfR4KEtsKx5fFkeSvRxZYuNlULGPuvGaaCaQbr
Ptd0voLeDe8KMaFGwxNPt43XRDKQwI/rwt47QFalhpME/yRZLnK86WHQGoZOjcSR7eG18mgyX8te
j87X/+xh3M/OSILQ/x4WlScvzhzNHn4YAf5cXzsXbDYJtsI7eYYKflLz+1AXj4Cyxj3o9XVzOB2/
upIIL+ypQ6NmWWkkIv7k9oYf5Xg/rRsEOgqJO2S2TilTZiuICBiqOvksrO8ZaiibCQJqmom/MPBj
KNexSEfNA8z1LI4Evz2j1aYD+hFOKfVqS04Nj5bb/XNzJMIJSz6ADgkG4o6698ioWwaETRS7Hxa1
tQLWH4rq3LbWNAKxCzpWwK3CUIgBJy6H+BMG0F8ThB9tTcSKyH2F6wH0giAOLY3sd4OXDGfDMXkq
DILi9uORmIoa2pKWIpKCz5fvTikmfgsY92nKu+Flv05DIIYQFr5rLp1cpApG3vOHr9vR8ioHdB29
UtVh+/tIWDzCppjpprmoVUkP31zhCC6CBObgq7TTh0F0EGxBTp2DDCUXGW2GCuZsy9TbTsAIUSTI
OF6lESWm+mEfD7lO/4uPndkaDvPpDYoLp96S8PsPUqA5HqA8xsdpTSe1QN8VKznYX1ApKclIJTUF
6U2VqjY5CnajQROHDmtmH+aCjpUewU/juLg8EC+kqK7TuZ+fO5lGm8sbvceq/64R93n3ay0FpWXd
OmG8es66L1gfwfidcEQd8CNp4ZY9AwRDgIR3mYK2Y37vu6OsolHNedHeJjF9tlKg2dwMNgL1PZUS
FlkX10xM6IazodpUMCaDYMFdSVSmz4P4roCunJLaK1ddhiTO8eHZtnw7AMmzk+PWeUV2U4I++Keg
bTGpgnnQT96MEtrEB9hEqft7zXUD0tbxKj4x0U9Vmct3iHgJbfiK5ON5cNoJrMV0kx0pTJTKiy9S
ZX4ypcZTuX+2/Vd1d5nf8nopwpX6urY1eebEbuus0Az83etIGomTyxlQH12LFEQiWVUAU88Vh6fE
wShYA20W5Re9EEb+fBkpUh1jCp0og2EQ8+1Ot4CytN3ZWtcnsKe9geMZEmedWRwU9jKYoir1a5ds
n2YGv4f4715owq+dVg1D3QGXCRHSf1u6hdTw9SzhkxPIepoY00Xoz6wLj9WRrkP8bBqspPaju8ar
rcM2YB2DxLetBHRzku3wiuqbQ3ZD4lBBfCXndeGnYiNNE+PrgVARAibycxjFY/R8T1K515ak/ANb
qIR6W9K0owCOUc5pOGNgbfTt4HVODqMLBgrp8Mu7c7b72FlVn5ji5hTxKCzZREp4z7bc50P9lQkE
A9g9B7GFYoYAGHq7CkNWiKx1wNVg20BUFsSCvyHMpWX2Parjc3kixN4r1AQ81Fe3qHK96l8kXrbh
4mobt23rQkF57SVOCivtkCgSCbjUd+x33BcpIlsKK6jLpd2W9ZFGmDY4ASu04MR33gJ+BIrk51o9
fcyHaMYJGYlLISUhR2YrWkOL+eIIuPRTgB2JVJKxpiJihOyMiNo9Fc9glODC8A4/7HA61gbbDGWe
dkBCCSOKju4WrcM1qem5wwGumY4emRKPSiE1SSb/Qki4CSUQHrq+RS278xXtE8n6+VjXfvJlQCoE
9Ci1kvqVYcENC2eG4U5ccOe/FTwPaIWDyiJv7XrZY8buQ2SQeahY7q9kOCplEJk3lOeYKdVHrH0i
BjGoHEk99LYFVwQ3ZdZt9DqkXxzRNf3M1czv77SB5t82NQxvXC1AiygfafplliHCwnpbQVy1MecX
dQ/2tiyWw0P49vLMA7QDDliPdu8JVLpTZCEhOdA8fjm6+IKZdpDPuyFEJBJ80EPB0AzUwQVntYWE
3EoXvwF3DjJLsHE4BogEDR+JSbg1LpFD460ysPBExNN+S4Bx1Zrez0NrhCCDSjr2xS4pLquOVg9j
kKYkTyKwotddgbAmupvoIs8jKZgRpaqkNVMwawS1rL0FycH1I+iDyWYGJUf4rG6XFMcfwFLCIf6o
FNUBxNT3+tXCjyd+DoDh1xGEwnHh8dhGujz/SwhfZweJQipWEJlUHAh8hMQAUEO9GJD5KanSUvue
Qzw/7hPe/GC6RMmfGNSGYMCpiEVSs4YMYMOkrkRX/5e5t26zwUC7gca9Nbhzz1UkfYH79GOO9KU0
WeYv77OYb6/GQGHwA+pcfwLON/hjtlwR9DWY4HiZ1Al8yeKuP6xBkaqPzZJ0MgCULSyX/uWKuA/U
TQMyemZqnIIdZlw+4BbYtYKlExTCh9TTB1DKGGTPN3TqeBGMZ0FzfkGtANlK7z1vuWDyPIAVYyIV
ylGe8oo4uW9J92ZMcCSNZvIuAJiDmguV7YCLnHryjAG90TcV5Kv1kPUGbGwvlm5TVvtp+t3SBBw+
PLz/HK0LAkj5fXvKvK8yvuKiiBtmICEV+glo8JQrVPdef0eXVohL22bLAXoA/JhzJXSy8WLVvBAg
C8HSqmGIbrSm7oo7Tu0ZY5T3fUlsc4bHRGI1Y4bUz9AzUXrqNNEmMvOBafaTXWPO+9CkdV++uC5v
8Fqo9h0rCtBxSRltMkqT1B34X4lAcaLAz6m5DH/6jueopkTnk1X9POd1nlQnieG0/oc1lTuZKP79
ZTlqpvXxfCU1LvBzMHUx4vUGpikceivJQUlZIO4pLcdOruxqtHOWU6bcO4fNeXBc2pWEjmrjd5+H
worq4ITahf0jwwQl1dDCaa5GvYDsy4TikDy75wZqKuEzvP0l841Ifyb0H1kEfQ2IlkyZ9o/dLjCf
HharJ0LpacNoNzm42RMphmHPtOSAcV2kdbQVmf94qIM7vbeGhunf2TSEqLC6epRS+TrXjUXZLfaY
3Mr+Gl11+bDsoxLwndtHy6Vrz2xMbtdFxgLdzS1+m/iDF409FiQdLapsiHzzuhLwyh/S544G9r7O
J/D9EzezML2eBcsKtOu1xvhKjCpb9VPx9xNaW4MtdCvL8CyrfIpiJLQK1KfYpkhInlLSYFdns0ib
WTcn6yCxGB6euSJJXD9HWPWvDwzTPV4cVTrPZtADC7FaLB6ngItjz+JPRY1TYuihowOzGvslmzdS
enBstJkNK/tLeTiHMH1TB+GY/uSmgv3wX/g46OMR+sNut0dZC+g+etHvtC7ksVYpusIhRIdVcXNX
h1V5DQ/+vBH4H2FgaG+mk7Ws0V5Z4mNsKJuVn8/wIenQZ2UisZ3ZEIqDjmD9X6m8bzTGckuez4n3
UogylCooeG0z5ZervMwtbf6rVmq/rVP6M8u2a/gbM4mjDrB6CzYXKYL2DFoBzp5JMZ8DM1O71ORG
+xiEQC4FzEzSlcVxMqLz8Yy5x9OVze36rVexaFtr+5lC5TowhiId3eyHNER3tUjSEAk+AseoAfE2
LkognPHmevfSr2AS0wB3hLfw0ZgkkDy742K/3AJA2SK56+2SZrwiqOwDrDI57BIGggsB32DLGTX3
yMvzrSJI70oU5Nt4zU4c7s5tEVHo+pkxF1r02QwJ9nuNu6zPoiEpckV+eFkd3nmNonjQqKgezJCp
JKgCQWsrN8nFpKWcSauqKriXeIPXGhP2aC0KHi5Re+S2BZmeOLfWkzycWPvEAsVPdy8iSTEzjiKV
M/jF+dQkj3bLX4VbemwCT3dknqrjKLCZ12vXjbJGrMSZllMlrBxp/ovoqQEg+HVllUrqBonUP3+t
imC3PnnIfPWKh0+oCA4v9Q/CfhN+FRW5ckZT8qD7iHMgqg+2wEtcYO923WjS5yZjRRtzn6qb0aIm
pA+CK6/1Lc9mJzzQLLQXhkVfBteMqp49nZCm+Cu5NC4KJ1Er1G/15l8gBtSJzYPVPeYfW9gk++kT
Vp4wFoVb0BSenlL4WFb3tix5+14uUSFZNUm1YO5amoT2iv2L76ug9e1xehkFV26nQg7hLNLB1DTj
n83JGDg5R3IySR8ousllg9wTM4mFcYOz2gt3cfvhHANvi4gtgbqfUkFakFVxsSEcbfiOts/kZ1aR
wLWul7pSRY9De70wzUPyggo554zp7pGPUQ/n/hwOVCJCgxgwTWVDlOKqEqjiqZs5fSWcc0FAYIgg
rq5Cla8w4aQAOsYGhk0gaPJyoX/pKtlxyINPAfKYT2KhVadx2iMSfbWAJIG3yZD3apZUVs9G/lyA
zIQJWw7YEWwRMajs+ONSlU9HZKzkJ0MhPqw/3GaOShdtHViZDTAlRh2IZv6/eGoEza3YrGV0QYyW
vaGCWBQykFQwObtU/SqzqnRE6SlySroe9dTG3VJtvFT37nNGEuqLdTAuRYT5R0TKzoSv+tJvMc1s
pDktCoOQGShJrs0bANS7/m5XnzyWvOLbzHMKUm6LY4eqNN0j/IXHA8/PULT2k6LhArSbFiu+IRq7
fDrAgId5sNOI6yD79r0FATAbiRYpYJu3IhzDnPNWnJvdOTXA4ZyzspKBZw8DEDsY4xrhE//yPI+m
DNY0wLHy8uog3Qf8sO+YB4INOPE7wwzZOFvlYhHFimeoGEBKmV6RFf0JHmtFMbPQRJULJV+t9SZY
eOhquah2k8pUPxZ4DZ7oTytWjc503/6qwTIH8BPtAWTrecXAj4RdMSGnSpkyJhkeTHsr1qTJFa8p
V0ObD451ZG5zAEE0ZsfsPS8XZtkmzjva0XlbvNjqYBwpwII6nnSKvOIdzcYeAJS/p5iIt37C+fDr
xHKIC+KGojS3pBGZUh+e+DGJ5NcnY2f6jDrxrrny0kIyeuHdRzG9HsigcP+rakp8hyxogn7hJqAj
L3SgxWQTrD46mrnuV4WuuLEINkS2R2KEHEq4eAs9F9LifvzMdZ9yL/PaKSjQiqUh3wkMOFRv0VJ+
fUUSiUNsaoQC7oV7rGEOq10TrnMRrR1WH9cnQOXo3/LbMgN7MpOI75nX0x12Sigrl3+2D+g8A3oB
hg3MCkObiy3Wh5BmxQlPSFH5idr1r/6+Ud+PuYyy3rtQH0CMGz8FJgM4OHA9tr2foXkb6deXQyts
fs6nxwS8Lz+STRvNK4VChKQrUUHq5jP3cW+r10qsI3j/zK7uBMazGrUecCCmlrCCcQfb7xIAtQN5
ohtXhaQJ3HIKtYZheCMzbITPHwwQZjcm2AlN9bwLuIXu8yWb1gA0UYUeOSZFK6Y2ItOB23osqFMb
Rog+Xel6cEllR/4KscG4V2IAQq02ptKbjLP/s7TSmstwjNzx7S2Od9vcCB1mPX7n5cfPbPR1fRqx
B4AhNyj4qyERHYn3zrxcgNc1f07I68j0C44mvTgUzzkCEDaAKsmxzEjSRhacsTWBmr1u/8VFCNKv
qAajAOrIc0AOUvZBYjm6kqCfuRL8uL65I/DMFmzmzZZ2R7JJg7PjvlZX3EYCBM8+Ur0qdV+I81t8
gcPcZr4/idGkdfOBq/gJDur0wy61ehui9G4LRhsP/59gmB5TbbQ/wGxrTGh2+IH/P9MFU/RfG5Gs
NeikOpM7g1Z9tV+uGx7GXKePe5Uf4vH/eXWWjTQWJKGgXIlO/udHvxb2212gLIEPpZoBxmWOI06e
xSn4BBMvHAbFm9aIqj5jnUzZ9u4aF4MqW/0/4PH+NSwUz/zzWwLvuqkxkNcAYt/cauZUnhQus8sN
sWUGm4D8SqGTwh498AnVf22nrX17aLVXq4z81ceDE/f3Orxeg+IZFzy1Ru5MPwVqiiEb2bw0Imdx
1hTDNQatJ87djemN00xSybClxBm6Q8U3D7j9UV9SM4I5KiyhSzLDG1N/bzfC4CifPzpPL4jus3j8
0oBdG7b4TrY3Q9+rqtRPlRvxYOP7DOqdWJ7ZH2+wPLK6sPDLTI6GTtnm84C8jCX1yj0kjIsXHJWi
86Rlxz+UMqHEbZQtOKbJGCK0tBBlqeK3h/v2hdepHTbCKM2cnyFc8LQFrpOkkhrDtk0EABHyNFqH
sIkHrmTmjwmjuz0NoVS8mz5A6NkGVUeVUGwngt890dK/GjfhcD8DLdtCA01NAnD18QCd7gtkXVDz
ukELFayystuMnVweYynhprR7KfjjZAv5xmYqB4fcaewCUcFsjWxfE/HV5fcNA1tmAYRis8bxIDaI
yD70OmcLMN6JyZTANU8rNQ+HNKKmu86v0KDTTiqB8W+Hc2w7Gi89kw6wUOW4uUGUSvaZsmgrGTpT
x3CvdT1kDQ0OTuK53D3oOHkmYF+yJkP/SyxlbA0wYevMkt+e1h2b+hTWyxJLz8p0EbzKxURhSYCq
HH8u0B62rfyr1QFLsaFL3ptL1hOATXPBYr2M1c/t28rcYVSeHF/hY4WGW14zum4tgipRRQovxPWC
7R6AmJt0E7R1oPjYaxaLJM46FpjSleYeCIWZrpvmB/A+VQJII4x3IYFXMa1hl615bGgi79M5IuZQ
7q1M6t6bHy8H7OxKb1pVELKJA6YKL1ICWVsb8WWM/3aPHPV/IaJ8A9JrYQU9vAWpg50diwhw3Dhj
xCWeso3M/+RbVde4Av6PrdY9eQTReJ+Vj27j4QrM4ZdVE42KEgp93nw8IR1GQa+3TRfkEPlAdINg
yKvu6lLVKqIHGTS1V5M2QLi1BOHiCxiCvuhRayVhM7xQy/3C6WVXZ/5JY72QTayFqxj4/9sDminH
NzOMFJW61QtPg9BqDClvMRIQ1I2J4rAt8r35HARA80V4xqx9Lzw9YNQVYihcnHiPocsjTrUBW0VK
g/AORBK9/2bb1evhHJBYLG1pseZlNYbJF2QAfnRwCVDP8TaNwIARKBj8by+xB3iRuAAHzkgmOfJ4
TQlEjixdErnxBv00Hc2THNzFLyLye9jdS94V9Ele1mPvTMY8yPo4oTE7+/t3SFIgWMWRyCZz1mDn
4Ts5Og372l7cOZQqjOht+/n2sme9gCMkjlE8XbfZuOr4HlpxLhylTSUOE5hIUziEmxn3deCcdsPB
IeGt9w1XhBt4p55QO9a0Y4m3TPiufbW+dInqsdM2UFvt2bysfMidwuip7MUqMp0iTFmT9oUrdW2s
xfJfyDLAuv3zgV2y7FcnNg3Nd2vjDFUshRJ6J82PaVIEeoFI4Ug6dFF++R1BUQUyuPU8FV19ierC
Di+VVsjuHU1fi1iI2nRJObvl4j2qnKPSnRFv1oWwrMPW/lPpu7Jdf1x14cPLUA2hWdTBOOJPH1My
0RdXtThyDgXrMtbebEYow6cpP9r3KLoUBB+woQu5alCG2IUrtKeCWJtL7WyD7eNwbdoFRDkGH8cN
45FCACwmRvkQsVVCePKrbQijIRtk8koO7Hc78vusRifK399Ry351A8AG9AAsLsyvBSC8VjbmtdIh
PtJvOEsS3L94Hri3HQV8Rrdlx6zwO6hzO8eagKto+Suh9d/htFWeixUHAnzuAMFuti5rMUBDXFzg
Gjj47gkwxLUnFiyFTEOsJeAlytybjaUrVzctN7IaDvTeef9Sy05wKA+Q/rYDnnYE8PlOXupiTKAX
uzQ1qrCgLcFrXqAZWk49BHxPj+ful5el1/N6fprObzXbMr5KKLbs3Z4KCgkGy57hpblGMSueO2o8
tI8NfSxpBwoBdwUjOWjLZlAD4nnimvUNoBwLC3ie9K4xCYy6p+kEKzquE3LSAYKT6wSYvRIBSLIz
vuEBTSAUWvQ3cS/d4y08D0uFDtf7LZ1DrENecg96IXgxPRMJ4higmJ+BILOQG5PEmyZ7DyQra9J9
nLctghhowMSYgwLjlQ7mclI5oBGhJJiNObJf90VW6eav6ZopdgMMlmjr/OA4kwKlE60nhr/TcJir
C9EdQ7q+m3NRMWXuSP3QqYOM9vlI8pYxdP0Fd858Z75eAQGqWXAklyRCwfF5pnGWvJL2otqS9DNi
6XPoVa0PTkFTtjE12iy473VmM6wOGvHV9WcuOqU2wk36Ev1k78uNG2rFmUf5Ccj9Sx7uODbwgZEf
HgrpDfzqabOgeQKxd0xALS5AmeAinH9hLW7MqUkGIqSaPyV6UFi7sc2xQv6Sf/cVgRAtI94/DXQk
dpe5jdG2IhQNjmRAvR5YStchn/TokK4sdYCxJg+VrZhkj8ADqSbttIfiR4pjXRaocPQIXVnUONpA
s7c6TVJYtTTfs+iImNz1pLbG5wYVHx7fn7o0tRaufRwbATZb3OVEH2iwHR/9wQfXBa8Rh1CEHvms
MaCb3W7Kbp12S4Kjv56hFbSmfMOob8RMDGtqQa1KIo4hel4rZAhCeWniPn0/zahggDAjN64kCZjN
kABypPPBz9eljoYfMSv1A6wDgFiQ2O39zXBhclfgBHa6lseHnWxm7Fu0sjIB9hT74RjXZz/LsIUN
3BP0QyqE9HsmheZ9trnC8nOMB9ezHgSpjwq7D5wpflJasH/kDycfml+GoVSUdDRt+D8S0UKQObwx
7zYibTgXKlQxJCzWbLdsN2UmdYp3udVws6VMFl3aGY8P5AdsNKJ9sl2zYDXyOrfU8wZ3IFfbHbtg
TeurngnOU95OP6FyeRSjYWXKItFzO/Nr0CRZmMGjrHAnYbZvWwNZkHaFlX4dx5KFYbPUzvVgG/bu
7tZpZ8p3IulKELugXGCEmen2SZc+UmkExB4eryFgLhqWs2xGMk2dG4hVqYw/LDxul+OUDhCZzevc
BA0Zse9rOePhE7N3d3CIZ5m/V/nCashmTntLzFIJgIvkwfegRABV6u9+C/nhM7o/qM39uEeB+nqC
yM/kLnhHANqYEkkXKz7hYjEBk4TNgzDjUxk4z/FoK+gObVh7G9iAA6+REjpAklIvns/d3eDr2I9M
qA8lmJoRwXnj8ze0D8ukpVo8ak1v5nF3g56UCOQk/FJJRise792vG0M9BCCEL505J9RQW0xx0dwQ
H2FTAK06yZ8czePJOdGBoMHjbVg5epWcRQHun8F5XBLRkSbNImfmpBbEPI+pin/E5iJUXB3/mxVf
g0Z/1KVtLiBKpxG/NvF06mxsALfSRnNbL1dWEk/soe6/R1aVO4DR35fH+JB+dK8bE99aBed2zaxb
PWRwrRryRxjY4L2UOKkFIqrU6fkgwkkHZyGwNeIYsGgWqrUyXWuX3uh6Im4ur2MXsTnOydJMcti1
pcboUFie8b2SwA4pMo9ZZUFk0JACkMHaygrLsGBJibJ3sOWxMJiwoAEh2eQ7lF4lxLuivFDAMITu
lKX6fq9k44uYyDUqN2C3cwFNujTxjSi5UDC+TcqYv6wpkQGWRyJ612v00X9OadTYdS0S+ONJTYzX
+lOgIqYI8o80Y0Ok1OxuU9xF/CEgtqp1WyCcEWm8lUa4jFm+8nK+WGpZYswkO4EX70C6v/qQBpio
iyKpXx7GNQ+E7C27PUj5IWTenEH4BGHb6K3MC4shBhYNSPjjiONjajSlQbeYaZGuZIvx8CiVnlqv
UDabHk1eiv+K6lcUtkPZsbs/UsKCzo78XErDGgAvmIAqvnVB0qiFwFThWDsheIDuQeH+iWqXIRTI
57xZW3tg77YGLboJgz07uvu6lYJdRw/pbETwISuqXOjtq5rMMQ/M7Xr7OMVvDQy5TUc12fMeGKcH
knvRJukt/bJgD4RPzgYdjA2jgcg6Qe56ZibovDaa4Bt1FcQL3hJorxbknJ4CHdAubzNSmIv7RY4I
1gEhZz3RZhv3x4ZA+qXXxrf9Ty0eGuOGAbDjivIts9pxpvT+z3oy+x6bCzPzXq/TPcg4apPOkKsq
n5OlvRWSnsrV2BkcApULIXl0C/GaSX2z0NAg16QQSgocww/U0pt1VMJkxie2nS/AU31fhmp49IHK
1uJ3iCBPGQpxhq06x3uUDwrIPbhHldCl5iRd0wO8TIj1SaJsega0RrBR7nQSvGiKjS4j4ikBaUPI
kxGUXIQeEiQkuMnDgnP53GoUGmGuoWVuZUGKNqp5MovBOgYhHbB+QCSIdOnD4gwjlMV72bj7cfwB
+x3csEPQgtyBDPo6iLzwwrCWPU0K7fc1VunCyCh6t5jCgIQGmOmrq13qa/X/G3ckPsvXq/Dv/+s0
cvD3yhtbvOH41LagzeoJgqvyQPfBCieIiXvaMUeopzs3NVoLrGG8wzMdcdDFZxbHuj5SFlO8aMH7
xxzSlqgtZdJNnJxL8qar0zz91pxduLYKidNFiOF3L1rRBJKdXCqDd412bvonaceZJc3b0Mvtij40
5UtB0pkCem5FpeKulvuGRQmi/4796QnNyAnZVy2beAzEQaqeuFwZbEUFoL7plhjAyPCcCk0CBi0p
dZlWqWhplIZlvrw0fvIW8XJrU8Ma/+kxJQwDm6aW9dRg1ZPomgLWk0brDjEazc+gyhXgLks3MOSh
pc1COHnkARlFXLWCWTiGgJ2XpOcslr9Z5wnSM7FIii9AhSh302imEi7XCf8vSWOOIhrLVjVJTwL/
uX1+Vyp11m8NlOZ7CA5JBRRTJMulSNNMYzY7X9s4w7IMpjDE0Yt97zZl/C5uBnNhQhYkWbcHm+LE
Ld/UIJasYs2l1Ef51EatkfX91U2SHjSxJPgLXGfi1MN5463TPn7ZNCrYGQVZkrRr7wkJ+OoJd1/n
VO8eHDUv9SL1TZcDGs1eQEeXRt2KDyE7zquOxWWyc0ntFicaaZPJVaN90L26WGJGuRLW/DXfeie0
oOrN70Z973lEHSW42ZHRUEVc7LLAU2+iIGHVQzOlJV5dTa+hgKQOWkTLofyeo17OECXSLPD9Lr+W
/L2Obyp+AA+ToVe/+NV0+9utPGDKiN8dyGE+mVoNMvnZi6bNFkLOJK6lpUVhz7Q/9wahdjxLn19Z
h5QbrDXSaZjKlwopXixCn+gqUf3xf0/ZafQmzU8g//eFAWTS4UYqvBVzMHaQm1hE9kGe93nSgdzj
9RjdspQ9DnHVJsnzrumeFnjDNuHJkZSUhQT4LgZrzLl9zYAWlU50nTKAW76+t2HTsOhQQb8sONfF
8dbBmD24Md0ZAQw++VKmNauDlV0I1DLldGG9Rs8ywR7cE499zOp/9GNYJePgZBdHQGYj9b16o+oF
ZMmHtws535tpaW8S+l5MQdSE+T144kWhpiac0dLDtOEcuyg0nVeCGFC9ZHSqFYcoJkdtIJCyiIDd
iLex5gQc93GEVGgkSHbpEUiAL8p8pvoZ1yW/7nGQ9/WktPB0rGWv/RtAPwRlpu0LZbGWYu15BYnd
c+S+d/bg7nhBrU5t2pIup2Lvo+z5iJqm06rudWfEi+9VLFzd6E9YdSNaOpyro8PccSw2VYIGcEjl
crXFeufx20kX/o9bhgPpUXtIdj0xPS6KlOcpamKWUtL7oU0R6XPx9Qg6BXcUC1MeLWLHS06eiyP/
FfzQBtwK/cNeq3pY5lDlAvCIc6UwA8l+B3fYjsKn5IyEbragWJPiRPB+1V3K22EOA9JaqkVgQO8D
xoEW2Zp532p3wjgdg/t/Cl/S05ZYMI4s8UBOrAfhNzJiT0UD5LYkvmq66dGQRiHZ9QoD73yPJPMv
bSZawY+NbpeF6mwwgKgyOQ+UUbgCZ1Fm1dNPfm1Vv/wtEd1K8x6gn+h42GKq4TBsv+dVtMu8TzEq
rb/Ej2Lx1fre1uvNaNVILxFbLl1gGx8220uno9AjSIwtYuBExvpFzu/XapxB9EgljugagQAn2pyW
VbHMPM/8vh6tWbzRobo7kr5FcGEd9X3ECxBuWTqzc46WzlqL55TGhIglPUY8hHF6LY6ADpFl7s21
Z9odP2Qrdg7mIzRS/QGbilSzenwaOwdeEspa63/vZmzykMWuhiZQUleOhtcw4aby64qwoE9Q/Nqb
9WeFMNb7MdGXMyK37Cfc+J6eY4ullnG+/b+mLCZ2CKbZb1riE18LZwRtKV7aJEF+w0mM55wvGqTi
znxmVM6aBskncRIc8GF38QdN9g9SMcFABrVGI9tvpMP3e9/EStcUH8+zShsD59FKlkllsYgJQ7Vb
aOp45kAimI1PfU2u3o+OeECvKY34X9pbt40j7ggAUgGsZclVSQ0i+vPSdhg5FE6X6Pjj4lu8mMx5
sZhOkBPeT7o9J2/6KiYHhl0CFxqlxUaMHv7l2baaAeX7YY/VbL/HFwA7zMIhi+2RTPBrpRVLKVYh
K6NblzE++lwr7XAzVN7SBONN1ECNz0QpmlVs2zxfShRWO261i5DFUNr/+BenxGKhBdxDu6fCC1uv
TqpI67P3l1trChqMT8Ig1fysUB8sbLlllW7derfnXy7BUscA8hachEGzuDbNh2CCGuYjP2SGivry
slYug/HT0l6Ix92jHq7fVVX+9mwwoond2ZozlH925zb+YuGdRSnvyD1YWmh0UNiRINhjrMWqcVT+
HspzY4co622hjHj45MJc5w4NirELYBZ72xMRoyktc6men4UUYsb2gqAo2N4fW+0zZa+h1Lpe45g8
R7zqtmZOyd3fvkfS3cMOBXaiKOvFUZ1o+sPYGWX1Hu64cTeKutHUJR7o1ke+ECvkN3l+Noc3gonK
l1bpzIN96Bi9rfhuw1fLyxTV0pdTZNP2UU8LRcwqzCRgRouyV4E0c5vdegNGvkRblz5wbi7d0ion
R1OYHR892HagXU3M2ApkDgChxdrw2teir5BlHI4icXpmTiPQNfwUBKoqSCYPbHAwkGMZwBS77Vjy
HNX/Rv8j2VD+6TMFbFYQfa1iNIF8xLnypawxLCrDr4fLTwnxGPXfRGtoR3ojtEkIdMrbGdD+BFfo
IhJM+wNBn/2URH58GsugAfI5GWADAdULgMc4lgKJhE0hTe226gS0PAo+X2AmATXFmDPZSlkRcuvB
2MEtcSQ+2oP3Q0PMISdZbCX07dE8NWnZVQyRz82CW+rqd2D2RNCb8yib7MbgHh3Iq7diBjLrNu1D
tBymZV6FSVmlTJH9KQhP+6wbOFAWUaVlaVuNteWhCe2OvC5lnlvdFcaCIhbUo66rZEk3x1hl5y+6
4OJF/1e2Xgb4OHIWcL0er2NWRWpIlqfrDeWXyDX5ZOPJwab2q7FyYbJS4fhrYsYCkuC0Gej8EMho
NM9ZVbBJfzWY6yFqL/bKd/SmXtTjYaMY2X1/UiOobluaBHTgQ0utZc0dkXVrqJGmGAYEPAzMOmdl
P5PpRccPoZu2OifuUBg0N6Mv0LzCuM6N9U1PFv4lDpR/JlMJ7Oolco+x8JoN+2CSHO3ikcNq8ykD
Fn7GSLt5GNk+wHVf++GcOCILy6saRfRFnOGC7McwHaSAeAS+VlKQmSVKrPXXzNH6K7ypkFV6TG9y
hUbUpCWmpSRb6XfDSo2J2dQDAVhe78CFzgLR6azwzAu8byQ5S8YjIEQhLaziwZ8yGAEjbGXj1LXq
w+7HWnzmiXnilTx85VuzpMtKQA7Xua4Q7pEEimvD8BPeAs+wWSFHtLJrS25E2XWVLj2NdTXT8QDW
UlrIPT/aTHGE5L5v2MkxV2K1ismVr11kiijCBwfOe/Vdboe2BEIjz9Zxvq2WIuNENQSI6is69mqw
1xlXIpLuORW/2ka4m3q/qEyRnDJJM9Khic6WeCSvZPiZ+UaApJLE0g6Raopqk9X//tFFSBRNtFSN
gSjTuRcWo/x4OvrkjbAcJNVg/cawiY2cAhR2VNeM7MB7zSvY/ANh6CTjqgb3QSDF+NX0eVLSX+ba
n+5+O9Psh+iHHKajf/BuHPdmcuYsyw5XUC1vsrUWRxTX8JpaJ1i4r9WTyNNoOzApCo3zEinQy5y8
HnUsTqJ0ji5sLFksMNugvtbVvw/AQ1yOEqwJ0owVxXmQ9WKS4JN7Qne0S16I3eYy+xpVxZ/972+F
VBib4UxzM0ChgRsRxvi5fg0p0VSw6WyEYo6Jbn7zl3sflWc1qtQOuf4uzwEy7qwq/1PCczp9idnj
rW7UnZ6PQbKJ39LPS+puVLUajRp3tiDPEgHLJUsLPQb5vPi86t2TFfCvZ3fYxbkn1PDcX+vJIhSI
j/3Wj+G4KCRW5O8vGAhXs6SBa9XW68U3fcPB0cZgz/tsmCkrgp1CmIbhhnn/x7N9hgqLyvguwBY9
Hq5c4IgbYqdNpfgSOurDzDvVIgXNd47GkieuoejGdwhbGgvhx+HkCwtrfxnAGvBCfeuEHKPLOPBn
Lvx/bzWsoPoHXFM/BD+0IczZo17em2TmvyHCZ3bo+jr1/D88jvtjfkQ9ugjA8tIQN2pgRyVFsMrV
ky9LipliByL4dP73PkqGCFBE7DzJd7hVIdoHdjeBcZDhi/o56pHCV1zUo4OmmFbv+ub0NR9ptq+R
SOXgETEpoQqTmag7S34x1EaoJDZ7n6lnCIqQHfTocCkuRiHyU+EcLktDGjewsJyCHOM5kld51h4H
iCU18skjFYDnnjmdoeBfEjMySJZWdewnnEKrVKFym0ues1Iwli51wHbADjXaz1wCgyYskpAtrt0A
VfBG/csno/WzmmIJIkYTHjquaCYJpeTe8aahzYWpHev9Fb/ZJFnoZZjSpd9faDsDpok3F0ur4ozw
alWgqNAncCDTuge8fQs0xGaSCJcnRA024fOHmZCCPkOYDjofnU4USnIUsu96v5Qa3ZjANHV1iF2k
fOfOmcp/h2Qi5gAf5JuegihtmOfz5VUGoxyt3I/qOgvK2hoikPrQPmD4Q+v8sYa9l1dUfSeDzQcB
But0aIGl0F9GdfWKP5HH2ijM/DSCNcRTMlFx61DTtDPORqPu1upnoz5Aj1HlrdPahUYlPLoBmrwe
4xLZHklCVf6jP0qfts1prHf2QjpIH2hSU/UA5gzXGvH1ri1UAR47YsAJDMNVGN4ZOFKyhCr4MEea
MgUxnAjKGMRaNerFNzG16IT8Lax5rQU1XNgqiQlJW5uAnkTvd4PE3F2u0DtmX6EyEE0Rpy6isdTh
7MwNbuCevTAb+uSh4SXHDw5o2h+bowoUxZQaAKqJSSftUlrV7PHrEQSBq0eI8wlM3vZVjWOI5JNt
13V+vzJ52Zo8HSFWd+bWk+SZkzAsW+YQgpUlZeM2FGZEJM17qg4+DzLUR8QRUxEuWc2ggObUkSxc
5K0IW2giIc5wwASIecCEFRLop4Q1BvyWuI3HllAFLMKB8YzZacr5adNIi/n7iCmgCOg9B/kea3ey
bFuOxhRCX43eOCmFDUkN2vw8m1O+BKGF1KsrgZVS5Aw8xrlGDhWSTjS2md8keIbbvjwLt5jm1Q/2
wpsNQjPB5dK7xbdVCUecqnFAM7qV7mi8+thRiPTSc4u/FEowLf0T4uRFSSd3RUoLK7w6+y/RE+vU
5ucv9FCKLzm1LOPsipG0FoD4r0SVPqZhXkLKwJZK57pVJeRyGWmm6hEQnk4qa2EOUZkqzQz9uZZe
rARC4YYbS8NyUhDps/S9Y4w4xLXDvcnoHGsLOLKK1REZZBrTfh1nwEukWgrFIpZ+iJRE3nBmB0m7
W8vMZjRT78Pxmwowio5xfatWRIu7CNC9nDiHjBLlGnXasd3LUoT6boYdHj3gzq4qvdRJgzYYlbhK
zKHVtZ9VxJE42yXKWFIdsvfT+R3qcafBPPlI/C/6SMEDzY2lWIDbtsh4biIJoFmLGDHzDuIkmOEs
ZyNCwZba2aR6KTwJIiYYpNIxCZACmZ7GCgk/PamWP0N0zJnoOqfHwnwXN7lICc/8z5eTZkg8AmAE
HoKFx1YkpWAtiUrwcCE+AxaMJogg2Pl4Rwgn9Vs9IIuoHe2ekjkyJH9gHhcjD2o4RmJKv/8YimX5
58kmlkjT1ApO/nKJIAAhZo79bEhFr2iJP/U1h/9VtchJKFivLWgvbmZFWnEvlMT5qVfptbtVSuIw
eTw6yz/g8LjodUPGJRfVEgWjqISglG3xoA+syhKZV/3nzYFFa3giIfExK6KxsPr+dWGVDX3IBPsP
E9qyN7saibrz3CWnDW7Lg5D+lltrYpj1b6WIS5OPVlDGpMtYVVdBQwKpU+yHfXFN+E1R7mYGvtk2
sIuC5wlQTVibLc2yesCddiWpWAIDz6xTtTqLV2r64d2wrf++EznYL5qFt78KvFORzwAF0IzbwB9s
KPY3rSLwsHY+KNAB5hnQGsWa6X4M3i7T1Zc0oFRlnUxo6J/CMqPCt4B65f5nhxZBHtoC8UYuayVI
OSMmare0VdUPQ/n5fU3qP171WJuE4lqHx1FxhAUg9qdz8h1aTOsY7gnXvoKYY9f6y3XUAJ4tmG8r
hWBcnQ/88aEc1KP51cndABjGd3nwttwUp+ouus8xZMlir90kjerNwuGUQZ8G/QDrYigBb3QpuHFY
Pr2mtrjyXt16HIMjh1V/F8ePXBJxkWd7X5Vslo2BMItsRv8yXesW4KmWQzgcQxL7M57iGRqOclcS
PY8GCRCbLcF5Zx9mORiU2gSzxOg2AVt2AQc0DCdg++vRlCK21lSPGgbhodegDysi1kWDwvmykHGh
smHRJEafl0XacuS1YykL3FiQnReNLzuFau7LAyjiqLqboCYR2yyE/RbBWiO5DYpcdyUSn579gN42
Mlh5YfNN4XgCmVkWeD1wAIt6f9KyWHYxUS0BI7tQGWdfvbKYCxGNola8h83OznXCY2ddO9g/LcQC
hZjmFghxNbIUcpyjpPZ+KOndPVEnojhohDzqwquS6xKIEc2kFWmpiuW/pELuutfI3AA+Ka2WUgrY
o0VHkoKokRi/BY/2DBYqWQU1Vh8Tf7MmtjGT1z4A3H55rgqzmKBy8azdKMbXvc1xcD+IPTlyLzFR
5UJz5Gdomzr+Nmv1T4AlVz8yYMjUPx7iaghg1Zdx27S9wrop3y2Jktu9zZVElu2J7AXiPEA6QIVz
ALSZcI6i4Djxdn460J7Tj+D/J5PNEl8DN2NqmNiVdQrPLMzJFn/RKyW/SPZZ/kHKboHsBkonjhs0
8aPJmDnh8Vl80FhMx3Y9PY9IbyQK+GJcIobtWNw6VC4vSUvi/uov5vWgjiQ8LxAxvxhlg1kkovo8
lwvm8MgvsVIqwneZrA20J7JcIKLdgyD3y/RcSZSwFrN4XlHQMkW1MANdvZEhnkjngT1Z1Rkw8R0i
JYfChfOCauU5/t2D9raOV0ZfvdULQiUrjczwayUsNrMy8ALRyY8lPzOTINOhmGH1ANlvtSbY7f6U
PPeKnN+aFkJY47H64tmqnDL5eX6PTGvBNSk6VS0ILzePUgaZJcUHiFctJQ3+bfE8ZYcMFm5FfywQ
FICMCJAECIMvt149IvyHXcVY9Ncv2qZ3VNudC1kXX2e0GoPY0fKxNY/PEw72a7uDastZxgQ5JgzC
EFaCIvBJq9YJGx9IRZ0nCHDy9nqvTZdav7KZbk03fe4h8rusqiS0PewaZkyYa6QcNyVPUv0L/Lle
DlGJd9eFNIDgWEDEBEb+FQaREDU9lzi3MInL8xbQEPTPlZ+rrCNzfCTeij4auwKhiIINhMbVsHAq
1bvJlBPK+Ibgi/SBhvwzJ3/33+zRK9X99g88Lj9Bjek+tv3togucuAdKtz6srdFBRlD+BPx7lFR/
vLm6kiR0baLYdbaGNnw7ySCGQ4Udwq+zLSKOV7DOq6WM9kNpvTtADMP0xOLTvGgY3xU81BXguSnv
XfiROqbeC9v2JAbUr4R7AocoXcp45U6OOrFzhz2Z0LfC6TpH6SMajlv9UIJlQq3vX6dgVZBGAQ2G
9IZXqydRLbuD0j35zlReZ8X00MygoXmeJah8QgsGzEbsLQWZ72rggk2UoZgutSRTapeDqeavCPhb
HtW0iwEcZiIh+ctHa2wygvi3NKzevQLXVRjEMZRZngqtZR2zcHOgu++eHfJ7PmBi/pcffJ6gvRwC
DMuEm3lLFbCN/kFWvQGXIbvZCqM9rZ0gSjVLhq9WcvxNv5kqusMXadU2moyOkxECmDJYA/jh55/9
DlYj6rSkZNpl+IfKrngZJ4WChorkveFaWdnXtvxH21jsL52Q0vMI6Bc8uLtTDqhEYiO7IwxxksMu
cnIRg3XYUabOxdAL0QIMBwVK5NYwrA4SX1jLbxz6DVUijA1zgcv8jmOJrKWkANOTelpu0k0DrtwS
ISLQQd6RDwiQ94ZeP+vs9T5MedIwh5zdgIndxDVbExjivP2qceulVvjax1ajPhVwAJy+M1sR64Us
++4o/8+aGtYRu40twpZAMYBLww9/D9Ghlif6smBR9x6FHVmeRHJ3hzNbJA2CVhDNLDC3PdXxkmHY
BWcWKufe/cjJ+pAh2AOm0pE0T2fRPWbtsuOo5m0sn9/PHvgIIvZ9xWOebTc7WlfRhESPe2s5tsyT
3vVYGYxH68nv5AWIGj57oraRRqU+5Fg377yMUVcj+3nThR+QbUIuCNpYR7NEKKV4unmzGmVItDOD
eZ7EiNHPqv4BlO0lv2h1T/R93PwsXTD6iba+ZpRxaYniF2WtquQW6DG/hclW7rGOvt4GlMPRK1cY
nVl8bv4TdBliyqQuvSfMQ4bw/U+KRMf2lnso20DEp6HmoCk0upj0Cs1EfgHUtBW8Eqrwws6hF/xD
VehxYY2ukx+ItBdMhkd8O5Ack/tsgu1jLraqn7a0R/vMWLyMpilvN0o4L+uW/VmZtBegE1LVT3HH
4AiV1bOik/82PQl5P2sbp4zf3hooywAoJbKUBOp73pOqTgGNTSm2edLnq6NQF3xH6wgibmqgcH3y
JYGCfd9+gQ8bpm9+S3RFRwKDynv0MSlYgvTjcSGvSPVV4yZGbXx+pxuWx6+7YV/NOQsYKbAlWMZL
4r+VRnB1bPFobrQWvleCVQpc+/bbVIxQZF0MxgE/pTZ4UxJ/0l8leVAxtCuFTsr9nikBK63ZgeiW
3HVoLl+2lEKumYO4EEtv0lDo3x+T2f/qG0YKHX805P66E7yGIyKF/8w5o3TcX3gT8PeJmJKYo8TN
6nJau9kCc56fbeIiozrxBOyAc+gpsWxm3DH9JxvpMUgDAgKjXfjTW8trt/ba84DjZq7raJDYvkT8
dFXnftrnE0bN40NEGhhZDQelra7rLjJ1tgc9GVzaCuF6i7oQLlEi8W+1qLhlq5yvKO+rns4D3XvE
vJbEpKZI8iJfSs7FoomWxx0FCTaHogBveMkSMQVo0pAumdsFMH9rXNFQMpKsxAznXDVFTkrJRSaa
i/JTKbkTFU+KTGLYYVER3xzhV5RuvDiNqf4+Prz2+GacyUyaPFnnXNSUtGjFHdJyzryvtExPoLy1
oPb7NWvOYViuLyaf6Z/+FiUaatrSi1EUnqoh/RJLwfyeVWQkedilYmV2xHBVxxcfdHHYLv93uhZ8
sNAsTHDi/PvNFnHzrk7D8mWtO0bKimLfxPUKiw2Hu7RVUnQWukx3xShds/VFmRgVPXqOSBNYp6aW
NEkqEGMLxvILL7YeYEkZD/3QLSNG5rXeQLS+kvzU0boZgTwtbzSfPacMOkC7ng9cyB7UNw9iPF4B
WVKlp/K1xghdNwey2Krfjt+KLEqoZ6gFBMudsfNH5xEVBlD9MAsa2wMpSJBq0jT+dlTeYEPI7U3v
oIGIRO3yYSi60mpqwxMG5a89uH5qWJ14Dn+JgHRk/TaTqLJwPaV27L+DC6BeYPgwLS8T5W8/9o/3
IV+3/Ijt5r7roKnG2l20SIa2BS4/cTqqLT6/Q//yTSX5XlK//ItmBS16h1YcfLjc+u9pfEmd6M8E
xxn/TLesoTRtjGlUDX3DWsfYpZmPSjapUawTUAapQtX1kp1ruWfPnOJDvRDca/V2dYN8/dbPisTP
Hr5TmSRN/bEq0uFA8k1BToEDpZ064KRSY6uA99HFbF8Du+gBX8E4wOi274O76ffumYTZmoY3GMfT
VSZsnM21BEeYZVBX8ShtnN3xu6ggg8eUMJeMAMzcbpR4R+f8blhQanIc2rfQMHFT4COeryuSesdI
c3LYp9BMBrALbVc7CjTmWr2Xrg5fLlxl1jsTrYP7Gu0XUJjcnXxIEZuZZSeZjcSmnf6R2SIvuBx4
UN0L9mhrfEWqvaKXRFz9Y54NpGq4HOIzcGwvfesITkwS+Gt8TIujoqV9TkOFlu56rCVR/KNcP063
lh8ikfa+jzMyQyyZbPHDGG1d9WwaR/Sn9TswcXYTATzHpIBa6GyM7188/KdAOtVfm42UX2U7liwn
3j1iHnGsIIMbdKRpPdYphr8UVcmgT9JP+yYZ4JAOmnGLo+l4aslk6jxDcux8J16q9uUYRrq/p91F
mSG0BPJzq9GDGdwWS3sEyQfcFINS2Z+xAPJ1bvLCklXd7zHdLdLWRn88UHlD7BUroEFCIRNAwORk
CGsX4s42v53wSTtullu36bzbbH2kwlmk8LTL/bq7/piagMHycljf88gGRaQU45KLsmv3PYOJ+KuP
ktmKPdg1hxm2RZx68DvfJx3j/pWTyr+B15+b+XuiKNL5E8jrnNHaCv5R5pBlnUip8SR9pCzIf/xW
v33W5L6/iijqoyaZGoBUymM0HhtnOOO8im5qsopLRHcYDboTuC9AuPFg8DKW94v5K6NClNrnBVjM
pjGdyNxfw8BZqP+3WH3jhV84MkaHEAzUINR5tdaC5751QxtCtBat+b3wxr8TSeCuiv8RafJ6Ztkj
ywBwdgtPif6PlwgjmAa1gELg9Rb8y5Pgb1BVDzVMfxBBwNcxKKRhBTucqy/GSsjWppS/csuJyAB6
P8G5yDLbvoY8wLVcnbDqMuZsc2YVztMU8sqPrs62RU5xJsYAZ5Xx1L4PCq0kcjLzt8mSps9KNTZc
vtphCTjLg3+IYNK5/MqW+UlcxSAwV5rejFrTN468uosAPzpD9YJc06VHKOFgMlocv65u7BDPeMs0
WoZhSV2xGLPs4m80ZgkQzAJykrsKaIOeIW2kqI6UGvG5Nqbvo2lvC0Gc0r+vV/oDZZnt4H3nRcqi
s6H2MpyXfJqC624hS3Evc5HAjs1nMue9HmCaU5Vmzb65kMXIYjmZv83g6WrKbo5yMV7PuEhhcB1i
vVnHJiWWDRHebZx7kBnzGzHNRvkHnomR8UIxoX4OGZN8BhSzrRzuVFcrS4UIY8NhjNz0Oqkm73Mi
4mb9DiZ+lieT5nRtG2776WPwPyuI6A0fvYAq1OuAjDSuKMIZBGCy+KlQEP7Vkhp8MpC4VlzYxqZs
l9hyGv1j/gjl1aM39oVjkzvPW04wNAlxpVcd+PYtjxJM+o54kTm8KOC6LHyyZ/e9WoVakWbPWLAc
DBuqijoUl7UPrLNEUNORhfflDnZHLoy4wGkr+uF6HVVVSmAAkSvySf4bSo0X+36Zq4ZZrVvWf+Xc
ISHU6ObRgGdckYranB1csD1DDX+sPu2ujVLsIvBuTN2pMDi0AzCscL5XE6WISdex0hjGD4XBJe5h
zs8j3Po0wzpaagroRh8BGJySd795EELjsxFKJx7KEwnYQfs8WWktX5GFxazOdFV1frRRB3Af5tN4
5QSAldV9DZyl9KJ2vAQmPYI+9W60hNTKXJm0i9RTObqruPhxoh0DY116+h6G8fVHZwEwxH/1Dec6
E9L2h6kJj0OpkSiM1ILM7btYeIe8x6kCYLfikLauQgjLRMSrGm0roqOqd3Dt178OH3fxj1o54twH
qp6h/hbyQp/O7JgfXbpukTl9Nd0AEihr/91yI94vG3NMRf6o8N3NKH6QNOJIwjhRxfOoQ2CBTk2c
7WDi4TSzSzAFguhq/EixjwJ8B+ZhJMWDEZiQVcnUOYkq3YgTM9K5+oJK0gtHwAu5TzVYvR7B1c6X
Pz29bWSYegludNCtE+q9kp84e6ZEW2LsKwNxOCpDaIP89umT/MyZw3lshvZ5mc7zsrkQ0+qEq4s5
Dfrz2cHJB/FJYmbnOh3wIP17Cf/eUGwEKFrRdsr/YRS0k02hhkimoY22sbyMN3T3W41HXpsSq2LD
UfULochmbeGqhBRF6xOUicoUqf13W0NC4H+8BE3yubFjVrTtsWP4LQdbS46j06tfjV/s51JeRLK5
TmF59SdHtvDcF4/6l1JXN8O5yyKrbFZ11GkIC0dWuVg8nQHntdEcvobmp9Fd69QSPiZUf6E38PNz
EqUzTwl0qiEQWEj9itZesqkRkBorgbayl6wps8Jk87mvS+acZNfoK5HZYUO2kw507XV3SAQL7kD5
EC7jQSoLcXH1NDS161yaWsjTyAqaiXwshgUrUpsvdUKO/nlQ5IErGLt5rRyIXnmqZa2ymzokBqmP
o+TcwnZoPI6Bjm+b132t0OXF3UPoxaTwj4ss2dWtmfG/9resQ6ffEYMaljzFHKEp7Mx90XRzJwiX
yYbB6T7rX7zw0xL2d5t74s2qBDc9W2sskDBO9KYU95Ulz1gdZco7KxuCgdQB19zw770TKi0FRpZO
3/J7qvjmpk7MKG8ysu833iMcFo/8io/e+PlSjOgVPawqChicWLQIey7tjJ+xPsqlhayajZ1AdKG/
xAHbxvJ1Xv1997V8TBT6/ypWkoaartArfZNMVDbtxrlupw7ZLNxa7DAiyUO6HNtTQo8Ayeup+hHS
ZyR0deHdR0ZBHnXsI3DbmJT/mfGpgK+t7RUvfUFEec+bdKT+2p5OC2Qn1uLx5nVc+W3mE90Rn0Nx
jN93pHOKR7Algz0CJ4LJIzgjLKiGMiQjmqTJCBqsoyVKFL5JOf3ts57PNr290Kq3AUkdJYHDKMha
+iw7SaSz9EueoPaS4LCB7ckwBUTVf6v1/fOii54JwuNsV0dneZdmYOPk+XRgt4dQHuM3PmKbmY61
k/543Eo4u3u1MgNnsXWtXBkxPusfOfTdDw9wLVzfYclivkdi31WCi+2C+qUGKLudpLQqoiy/rJjS
MkLtFBLKdhPK5ZcSbcdTm+wlPezRYVDaf86XlJ+KSyjrDtIACqStQ7V2rfYPgDAZh1OJsxj42thd
W6j/dvdIoe3xNZhBMWp4EhJMHGyhjjYHVRi2qcILREbi1YW4iukTZgcegFB9d7ZJRKpAOp2jF+Ic
zPEmKYw1vMfkMoKXvo3ATan/uHfox3Fa5k3OIiaPTuFZwofPC9lVyzCIlZ3yO9tdlg59UkoavaEF
xyeJD1oBIlxqHVeNS3CHj7yQ2xI1KoZHq3QNQhmuFUHbsWeWl+xm4/mQJNbs1pqYYacr+sGnHHh2
PiQEulCKNHUWcwwNB2MVJFI1tI+IvCyBGFMoqcGBmI5UYTr5q8AmlsQfCo+8tAmxI8Lw7hlP2EsU
c9UnsRrrZkXoo6cAJOxZ/z2RoQC/DZ+TVX2IeEJ2IjkDfm3njGlqXju3U0jSX5/wp5c5Jmo2o/X+
0dp0EU+y7ml+ThrqREOhxJYSiIv3mobK4NL+UnSd7EWWFz1c7FgzYEUqzdq+R/hsVSxso8ZcyIve
mGXZLtvfRtnx+pUXB0G87Eekl7bhNHpMRZDM3fIYeZiLrt2a0D1I3Z0Q6xgSqO7dB/ouhgEVNbgY
wLXRWyGtTTbPFxXaMKg03p1lRAtJ9eJPhAOOEdVIeeGcW/z7EAAtn3KvJsWRyJExFGRQjTiKDE+H
l33Yb7f1ML5gIs0P4Kd62nYfLOKXfKCk4Z74dHhm3m4UWdjrUOcsH+K0++hvOqnF/7ICUwo8XNpB
LC8YYurdA15vmk5/qN9/gOotLTEktxaByi5S0Thw7Ac7Sp1+dLBOFcCTDkY5oZ3hnivSzz3iQPtM
/N7YkhBb8YCsd6VWGCF9IFCNoAlYyFrtwEV8TJ0NyILDVIbDOCeEzU9e9cCtLSzjToh1xBppU2Ro
OETF+nuJi63iTCpt8Rn7RQMoaiLmGZk2cT8OtxImru1J7plHTs1fQF//4W0Yzg9Dujsb/m+WBvWk
AVm6W5XNQeKxb4f4jJI3yZVTX70a0yhSqyNJ31Am8cVjJQT4khgkujQic3biWHDTQq4pQehZFuu7
+gs/xRNvhv7yaNoz0dnvxVUs60IzNj8RaDPJ9XGG432gcUygAVSv0hSizPnhyCKHUENMFZYCa5+Q
rTsBVIf6yNG3R1J7cf5c+CkVoHyvWZ7GcqaUzWoeHJc+xqQQ2YwF+F6PNbQ4rDE0u0tRh0ejrrdX
Y1qGIiPzHL2DpWYYpqt/zznzVZWQq1CMmNaJ6rpJsOpV7WFQ0Y9IyU85h+A6Vdxd1aPfTTQzzaju
BIhnMXY/UTtyOMxgKyixbLMuKlbFEl6oJBHwWZI47EF1WZcsenmYAaqqX36IovZeG1LTUE9qPzzf
dWSkHTH7leQeNOzg3QMc7oeT60VHe1oqysMndWGAN0UmH1LTahdm4kR6PqHbl7ogQfYP7MmuRpxL
J/QPXX6x6GnvNxQ+SkOYXLxFHZnJItfhvE68sRbPECy3vvX6fmg2X9m6hZj2eK0X2QhE63ZmlxhQ
NNguW/pKyx6PyTG1YDzPxcMJDNiKQoWnPmEGxueD/IFCDwOrQa8LZwzW6OLJ0IRahYVZFRNdnLTB
Y3/k0yFs1wbjXk1TqIDxFOhEr57qYJ6SP63PcKZ2tynM2eAH1hjYj2Bl/Bjo2nIaTHSqB/dllzzk
coY56L8/sD51ywfR9/Bwl/W+/I6u2EDGaRmHSaR/zCh+PdM6FXVcYrcHrpvApJGAJIHeiBhzCFgn
iZ+Ll+/BH2++cs+sBsLG5wFDaEyvMtYFnmr3TUPw2J8W6UL3fDyTX1N2Pn2U3MnlF+Vpz73CsxN3
5+6rBNaPUs7cyQI5LbXu7EqNysrsp5/XzNJcI3eLpBwsB6n1QKV6QSdVDWHO0NLe1jVHthr2FeL/
7t4OQqph8fz9qNylw5dhwyAJ0q8c+8dvY8QMxoGMqewaE0kype8yih2cgBkUJ7kEccaGEcPq5NVv
l4UhvYtr+MTntZMOaginLWKpWPpzJFioxHvBNJ/A6rTb0RWnAu4YL/vskqMtZsJKCaEx0OPFkLWG
BWqFlQvs/NCMoatQBqF4dWym/TdAMs9MkCU7BEc+mua6Xx973xevD6NkAcQ+7uyZF9eIb8FRNGUl
ty4qV4O79qu0Vm6aIcvAi4aJhg0fbLZKOhYXgtW9O6P3NiaIHdxlTpgOkKOIeboPt/R5inh8bg4Z
dnNmbsJKEj/1EejO0NRX+as4thp638Z4IH0sdNx7YyAl6GIrDrceoAm/Uq8PSIgEjig1aN+CtPfQ
qT63gC3LzpXy1sPHMzyR2qs334bPcb2H8LsJ9I9e5HV1+DONGpdL7g/2M+KsFaXDUrBW56fsKkJ1
N5shUb3cItq5/Ux6HxosewObucAMaiNU2Clo6uShscY5LtX2JjYuNQIgsSCnJCPbt8UnZyboODBC
H7VPx+hidHpSa0jgk5BQl8W7fNkANpZSPvzlnu1RhP8dx5Hx6C9+FO0x6iX6Oc1tSY76Z4gKddh+
za3CZ+yUxJ0pponq8tfPHPhOq6Fd30a7aH5ke+AKxkTTUe0gjdQh2ixi53Szfh8KfKh62iqO+dw1
dRhG918splIBa9spEfrNkOmZRmitW3/Z9HTnyHnSZqRJaoc4gQ/NX+8JdV0xSN4IzGycsgtO8IfZ
73w6EjCFbqoZ06sGHrYy9dBqsUyQr11bXiQ2pxW+/+RsCkqIjlHOI4v3tgAZBN+r0X23Nn81IjIe
glUsovinPS5Al6Sr/Un2qKTpSHioHglu6UIDK4b35xxkQHJBHO7KrBgZ07T7pIYsQQnUqcZkuNir
7lMJoG/Cnj6r/M2z3VY7/aftJRt7pkdUMCRoT92tdwcsVO5gZR4rXyU3lHnxdDslb5ZW9Wugpjvq
huIgX40rE9/JMoqj33A25hWqql7zxyhFs+4Z8NlEah/WQfHbn7+bg0qOuFLxvLkU/P+osdBGR2Dy
zvL1tSs+IEOAWfBV4ilp4W3RtdAdK6qG7D9BWdVjJIB7eJrUmZjFt68ssBAWfn2KWl1EcNAXJXxZ
N1GxBekhs9YVNsUcSFu8l1fwmxFvCsBTF273Y7gKWvRPkLSNJ/b/BfIQqEPf06M8wb5GYe6zjSHH
D54O+tJt/INHjugIzorCCVoMACpzHnhKUczvPeQ1xJV3prqRMZ3wLkupKRn+fP5VAeqaaqSNd6Lz
2tMqD5iu3pHgm2vd6Zxy3GkQViZLNME3lIizsdNz7gWwOX+Dk/wS+8WUk9aIsLdo2us7o6JHekLt
QahcFl531pBPyvhmrLGNm52Gvf2fc4wpR/vTE2DuFLch4iH0Jk2xWUsERdOrKGNVMw/6IYAB1C2g
5l8OvFF+9TzX2SOeYW1Z9966gDtusw8EnVXnAOfA2s+Rv0viKwHfiGKYa3w91jj+jugsh0FMYNcb
iIAI9uYmI1ozON+e4ShW+ZPym8JaHb+DY4+UriYQynznz4cP1hdN8EqXwKXTi9/TpRj+Zljo1dDR
bjNFXimenyJoqtorK8wZyEPAmfmHRRdfG4VToNTSADfa8yw1hCMszGB92e9mGPfqjBzkY84FPFIS
Q5q8+W0UW3U5dmlGRe9uCddMIxVaY3VGyTkY8enC632+po5p/vsphsY7VK3ShbiJQ8GafY7qyJ3R
Hb7sHvLkEKwIGvByPlhtpTjZPl7H7BbWXipYnkJpvfXkmYPYpgug796kiJmtqqRYUipxLoPbn3V0
n9rfUaoNNl2NToplu25stK2dUVM44xboFrsn566vksNB+LbkZ17tYuR0FcqqtQWetRh7JCjPfKdk
JIknR2SW1rEqHUoH9XaqhXni2z0HOFETQI1pXWovH3YMKqNmFqsNENw/nCiW2iZJv7l3YMgQlv/g
iZC9cZSbxWRJp5F9Cv89U83EpudQ45aLiUbODq1GAiW2/4xugkbMPk3ZNX61vneI7j6OwueDejP7
cKp28Jlk9wC/ZW6086fZDUyglf0gsacs9CPFCVGww86vjIhNYKTwJ1wwv09/qIAp7/wmOnBsoYjj
26RDtBAgvyxTiBQbKGTLYYgn0P8+Mg70EjFgftPz6aTdRb4GVxhRIJM6Am0IeoPW4ubJW3gZpyNd
fAHhnF0HiUmlUL8bFMlXr6ShLAHwWmHvIJx6gpcNG9yvQTn2hAEV2dmXxbx9RlWRkgE9g7Xny8Nr
+pLeQqHtITbfyTG1an6xN8hj7gjww+mVUGfKVkAEZwJ7SffhNbb8Rk9Uwind33+99A+J/L4KWcyc
Q22aHJ3hD+2yUVh5PfmUWqvY5VQbivflPGKnKGQCEmeBlWa4bgqA2LPjmJ9CMnSmn6Awtjr133VS
lxzNyxyEYxKJ6ITxoXbmVf51bCQag6DiIQy0nGLluPmxg54eL0QH/AvyTFbLlrRzan83QneEPhi9
7liSl6vG8gRSdDRCsHW69XnAKf59RnCw7TlLn5UUoGV1T13a6SCA998SRCqXMxx9cZp+Wzw0L7gc
mrAiH0xqy3y20s9ivzRwojy73pvnDCwKpAhrtrvYprhh9Dkh4K1o9O79ontWrXjl3qX31hU1hKhx
7kZGwVtkt9FFxzrUQLrLma0xf3Tkwx85Sp9xW3wl/gbU5lsLK2hG3T0LSgTVKxtHaMa29sdCPnyw
/+FY5Gq2+VP5d+IKqpuSFkBm2jQAdoBak2IU8Hc362gFOtfgKVvdQF1glWz7wl2ckppfUBluv7xH
JJ+3agCVRIOEinDwy9t4b4U73ukh7jW82+bw44H+R66fV4h6mFokoNctLqHW6Wt0HduCoBqsCEQi
wecNKbJDhBgYkVdcZjoQ0T1tX/VnioaafsabFcb/Sji56x+f13AQ14CGPwz4L9KtJeBwbMzE2dIF
nlBNJF56DMPNX52ucFkdQQ1YH+ODQOUTgZUzR/YPkor7RXaIBn/+JrhJSAfBBKV5/1H2FgayXEx3
iB5+Uc54bRtvmJjVtEwOFVNlsLzyP+ugA9FRvaTf8gI/jDVb7mtBycuwxKpsVS6minUjbwWFePjI
KedChwE2Sy/UdjxLO+5Xp4lMQ/NxhDNog8tDSHaWa/0SaYNz+Hz0eIN/dH3mBjQwq1/8WAeAVjO4
VWY2vMINxcWjp/ztnUoJCye5dXh7qYn+ykBUEsWblLi0M/LsFTEQm/2tDc/pp06R4TZm96KMXI+9
OQasAGDt/ZbhNqLXn6uhzFA5rxRrqHn9sROOdBjB+tph6WcQdT9+51KO86jRnKSObCMKxktGmnFp
jUS5FQ0b1McwwLWNykbjWL9lyn1kYQ58NnuAgDM6Ps7syNbriFoWTh1dmltrJtQCHtJWKRwDQafW
goXusacCEuyR3Jm/hFIw6hux0h92HPidr2GfaCCYL/wKicx48l/K/uq23g2aAvcTw44LWlvxGMcA
GAXek0MaQlFfZnozfkSViaQAPb9tQ/mC7O6gfJ6yYDUWqWtVF/vprJ2VWeWcEZ+O9EXURTszCBRp
rk/Q1eEw7LQ/DPj7FQ/784DbKL4duLTCWcng9Bv+7tiTvCW6Tol9/UmMyRSg9sIIA+o3F9Hb8aE0
b+Du6SmYk+zoH6+DBxRFNh4YZsZaz+NUTCZnEmQKx6cvODmrsWWlJCYJotQTRR1UsQaWBHM9D/fV
heE+wZBzqlgk41DZcIkMET7dfxitmvWp78PrGYLPfgAgk/p7pc5sGNVp8Q4b6ytrYVGn9t238Bn6
4Xs97wcBDQ9cE75VT6TVLVRM84Ox0ZErf8n4pAodBnATVZ0zLbzT0dGSYHPDocXuhvhrNSY2WNsN
8FghucGupdWQYwl4KRpKk1Gbult1nG8fxqnJBG/sKjrNfLRY8zAa6V5XIuvhib9X/rmK0igIsY4q
8MG4f7BG1O8CxqsFVNJms9GoiMMXcdQaTKV9FUMsQ496VTYd3+7Qs3/IGjwq7rErUdhCr0aoxIxo
u6TTpp1GpcYmVb0HQqxHoJ7W/aLgvVsAU0PpEg02sAB308nk4l2nWSL52lFsln5zYfbAydX7W9IJ
xgkZpyothWgFchBHEO7kjk5jro63ryQVQ08SmUj9Qi9yRU+iRst7d6Og5Ldyj7gNeeholP7X3QcH
smGBM+gQt/Wgi6f67BNgxSOj9ojAd4A/Y2NPygqv1avBO3cGHMe8zDA24FnKQOgneLfaI1FUzsn+
o/KzI85viM+Hd7rFzqsb71zOmeDA0kz69aNEnDQlokJOIBzuJToOYvK7npTvvkfR06a5sPl6FbKu
BcNcBR++TRp9z/vVwzRKvpLBZIeaMASSmMUc6Gx9ZBgUMXLAYXQAU77XtfHKhluFRCO1qLHE43BK
KGpdqLomdetV1oJicBuvuirQK6hRQeIdR9ce1uPxAdULh+lNTCD3T2jbd/+91f69x4MPG7cCTtjg
o14hYJmiTUeReAURustw3CgiIk5f5mfLKDsCdvwun/Ph6/KtNKDOnCzHOR5rfuPrCclm+YYg9L8a
qpoVec2E460irR35YjSstNerLZDaRarKoQlAkAC3hDd9GMXYiTvp7S/iVOn0/U074finC7EYIRyj
Gw7if7fa508f8gyt8Dvqr2oFStS8vPAvX9ZQEUjO2gSmqRcDdBkGZLeCUW0MIzn2qbsaIq0qTFg0
siqii4N1Hi6nEApIv8jpFI+1wtYa1N1mLgfMQKzSKWRlp34Vdmi0g1ZgGLdsTsUBdCzGYh7xOx8C
yO/2fJyvY74nhBI+fJAWxNSy5aAx1vhSE4NYgV+eSVnIOpJCBB67LxKxVzGdYzsqMTkQUoE5XVmC
5WDH3V6FUysd1QtBEvt3ll4u9mY5QeTNO53jBix4JprdhNwjjlLYPqspP9yYej6XAEBEWxjUp0OA
1pVhb7l9EGtE0NLyRikLaZExdfyQDgTJnpqyUynujORZLRyyRD3LP8c9zZndq1LV7atfjrJNWqtB
5317niAquHbeun34P5NdJzOo5RLWWWz8fTn3GsQ7Nzuv5t91wvAJx3h2QIO5cwTIJRxj3dftWx7+
DWrNRrFKV6AZpctf7+kknRkqLjeZUseT+G1bfGrgFPLIY+Vwrx1R+bmzEqd0TK51kJWeQvCH5pLf
XbOGORPxlh+eruHi24+/ybg3q5r2r2L/gbIqyd86JpC89Axw4UvlkcpGLzIyMlkHgU96ojsz1Ebr
01udwSy0/kcTprKhG7YAp7hksBnCvLH2dsKW2Q1Oa+XvzIYrzurvsomPCdKRpQkQsX8a+2CDPuU7
jsYuF+jGsBL/l7J+DRXiDXZXfO4tAG0fqP68722yIzh7fwmGsZqWdFTKPOMWyBwNXOxAGVDZ9ruj
WIf3h3MaT5nYIEb1pBpLAxPNIeVwZU5o7lRTxFLMLGVX8L5M7/vZr307ENRr2uaZRqtqkgrl03c6
uURCDLhgNJfv+IyhPoAnhcD2xjJVobLCUgQ9o7c/DpJn303SAXqh25iUM321V2Z06L/CD5HML4GQ
aA4cKqqpN/X8SSDdkHaaY9GWADDcEia8dqmDrMlwVWSpx+2aGRVY0VzuE2JlZ7kYclzbEhoVROse
zjAJJRup8xl/3nQUeBcBRvyu2pfPsYjQlZ1A8xnnSOxXGgq/7Ut9nl4snks13nVmnDvIjwjjVN5i
JY/u6k+EQr+Pp8OjVscBG4mTyCMoI/BdEcEKV91PdedwgLvo7MMIJAj1U2lJIEUPYtLR5TD0z9Sa
8vrAfW0m9MzbklW2UKEL7aiRuSTHsZrvYTTFyg1PzvSFzGeXuOJRHynIp5RqJyb8B5j0iolY4vqk
RgrK9QXDpIyqxr9h418fa4kXgG2SkSSg/6rW8yJblk4uMItq1EmTfjuYkGBdBHDZK1Q5j/h4StIy
I8Ig+HjIlGueuzyCVBVwZfaGEGnCjgMxWBPIKDbLyvxX5mP/1YL0Eo73xzt9566FQJn/ft6TIjEy
IiSw1V0kKyi24ddi+3skt0dJ27TG62DOfsmmrP8RE/A68qzwv/XKiMcDjE03QDMXQUWETt6jPQPX
YLpbeXfvG5nryw1hvMKh6m4jxf3wVC6HSw07sClGAK2MrRCcOXCUia+vn4m1FTOegn+BuNGYo98w
/bL1q1MH0VCT9nl6f42eC6soNUsB6UPUF8/hYzPGAjaaEDaQZzG7xrC2umVfml/YMWgN0FaOrr7F
MIIH4jOrMeFb6TjLX45rQ4SIMSPWckyC7CqIp0aKLXk38gLKdJpVJrqd6DJDeDpcWD6oGVrk/SuP
q4j3pxHhnBNr2gLC2DuIk6Rzo50spuTu31a8Rv6GLXKlIRBnVryxRe82Mks550VnxXwQCyBYhG/O
FA7d+KURUUnKUr2wVTC37I9A/R11TYijNB3DqWpbgNOlU95kOhMJtY5SS7QGW9bfHdBmMSnhTgB2
k37IcIPp3oRRbWwlFPxZNiYjAbN3ZNBHHaITe+dShPK6CiD3WgMH5Pttnb2Gg+yQEJU70u8qBDZX
RQkYvDxcAmaElpOzulBbh5uizNUVy7zg704RFkfEXQmlBbX4dJHHJgVZxtq8B5pqLbkefJ53Ni8W
e2vuUI9XWqyn/GXaP71T8qbwkz0LvIoUVVzWom80E+KegggJRcEyc4MpL5GcIhCUJ4N4NGUJldwG
49sbHvm+tIssGeR9rNiAgF/T12O5z4XQjNwmSqwq0RD5jX2NqqFJqzgyK+uWG30lq2YR1ieCC5Q2
g/ojhfZmvVKGdT+Z3WUIrAp/Z9mMU/jH9gzqwhVp9A+7j+zk2ctS5wfwv/vyVqQHgnl/pcJ6nzuB
kl1y+8A9P5KT0pLBbpOCiv+S712V4w3wDxWWpRWg3/4V7/IUAVOW8rlR/HzUM9DBf01JMOZ8yF0k
VsDQseWg57Ap7OgWgsr0T0XLr1BTXRt2Iyo9SMzaCW/RJxsQH/v5Tgt1zaGnZ1eJ00OqpkMWM+w1
MWxH60xNR6MWo3hVk6UDJOtvm1m0shWwDe8QBsrDlNTDseQ1hYjCDVWAMur7vXg2Ct7zJUwQLw1c
0L4o0kAJOOCBPYSKPnKAsHVj3xhAGZfM5lSuPOq0p0spTFImhHi9S0ED2Jwofr5TjQAONAoSEkuW
4gKbHuGznkufrR7XP1+HJyaFY9QsG1cq1Ar00Ch0edAlvoP1d51pguy0f1TB89rDM6KqvnsMhS5m
dJkqd7IdXNkcA/TrlKr37+RPAIIsLrBKAvpLC5BPDBBy9a9I0r8o4BSq1eZO+zqUQJbfX3r901T+
1EsbdTdBaFOWMiZvoMKW9UqPECt5eQNrZhDG1FybK1vgEboInC+n1XJzkpBoX2qZMx82b/cKfapE
V6Jkhj9VT8dqUQm6MD+Ze76SO9Ybr/3u0+lEar6pEEyd0TdHuV9HYQ2W7KZO4Ho6mr7xFBUwOx0D
lRaBtViOj0c8iZtVmXXz+523+Pb4eDUieZgXdBcCKyDuvxye2f3TkKyWm5tnbbowYISMLP6NDeh9
WEKw1inAi4FV6G3qQ9XvWe/WHgmnVumnQfIRaLAhvplRPNIuvFnW15lFtA1o3vTY/r6YMiRB/G88
kJTWfloCFz86vB2oJtt8n3DLjQp/7WUglz5YlgRRgiOYclR3dnUm7Wr7kMuJsUXpxXbdLTtLpVrm
T4lYE0IKT+7C4WH9ee3ms+LeWeNNBnczShQJqOIGaN8e4bQrfV15whi3NOSVOczz/4LrMMoEvBcc
QtwFIN/c2PgA0osT0rkVcxkj0CoCRxceOF4ne+ofDffc9RJ2YA7xUsHM/zyBssBrTVhiO/iDm2xD
Gb5v8n1xt9ZzuRmG5Gt+bbyqfDFbAwEV2Dh2UJZceiaGDBk5gAisTaEmmzr5FMn6RmgxXYV802RE
ykbQufPHKDdTYlGOXV/UGFuSKpCA2rOwLWpuauFWVSQfBnkBDvHxFkCWRVuHA3KQjUksLbPsD881
NnTFbwZzi1843/n6MtnpqxSqRFmc7ekH/iK3IuXipNb2/xQQhT7UW4oZ+AANzvt2o67x6PN9DEeU
7PA92Im6JIp1jz4Jj54o/ER7awYV12qegIIr0TFFA+tSrjja0Z40lOs+bSA5rFELxiuyczhvdKJN
FBbCfKnlVkQLblFcXt2YQy6bIbuLgG/EPH3A21V67lZ9ylpUpMf9RrhB+SrW93iRFTlkdyeN2M/P
d6BJADfkSUHVpZ1EM9zt9ZXKx9oGLkc7MzWOQZh6KepfXRDFYMEuhk/GZpBbsA+gxmorVhk46Gik
zOzQioU41wSFlnXSUMWsqAq+jxxbEI/HqtSeE9PErdFQgpX+82O1xoMWRoO3I1uCu23AVQBUqFdg
V2+1W7Ky7WN0EUczGerbsilAC28UpQXU89Dcfq2kCF82s/ZCcSw9vmBBJWhKJK16qjntcj6Jj77G
gV1F/gn17GVnzQTT8iC8jRQGnE3SKcBiM8FZw6JoWVsFKDFOqw3/VyrdHULXfOnPF8PtwCTb1XhO
u7LZXDs+F0MP9KMD2zwl832LZvB8QldK/A0VQhdRkibLQW7FxCl1Qv0+aTaw7C+0nlPrbqxzu1Uq
bPklJW9AcxNqUSEebJnd/PTq2BjmaXnsa0I6oG5T5t1R5SoDAf8/bRagOPrZHOmkQpP3brrqGkHc
d34wGFroH8pr7iDzBbnPi0yi8Mjhzsr8iIFzrz/7Knmo0+u7KgiQ7Sjih2vu/X/XCgKMl5DDXNf6
xKCeZSSXbqBtrEWU65d80M4XtxZ/rkawxbQwJwEN/K0wnWLeLIpaTNwt8Jsg6Hv97/q4YCV0CVPd
UmJ/nrfDi2dqx8Td+kCiKYLFEs3G29R9urqBB6iVaZlXNp0NFtHsTpwxdHow6nllcB+WqyaoSHhW
CKBnOreqZYX3j804bL4NPeKY+sPH0XfcJw84yB2DQmXWP4sGS35m8B8nC/pTp7D3EqSInw9q4tPN
Gt6fqFF3P959dn+VFU5KHYb/UmE9hTZlrpozWC3SwqWWDqgKiAruxk5cf4Sb7UrJbI64Fy9X8DSi
VRW35HHDmDBQgKcayIbDmomxx+j7X+8IrQ1fTIc5zEqlu/pEc3BmY8C3VzR2RXchx0tpcP/iz0F5
V/Krs0lVm2f7fxTrKTQBJ6KN+kiwug7md+S7K7CMFOe/nlx6bEk+CAlRdm+SGCiin856fGxbPbmp
u+0HHIRyePbPv+bdX7s1ak+lqAReD3Qm986M26Z3j9cjS4guqoUds+KNUrktUf3/VmKhre0C+kGh
zzn/EVSFtfi350vbn0faSss0dzhaygmen27zn8iNexh532e6VN/Ad4tmHzwL9fMMAUJe4qodkh6w
DEK4wH3TVGXcuFup+H2NhGp496aj9SlS8ajZsByXTa1Lzyo+n0nwtRACDPqKkye6tR1ypJqsyX5V
MYpUEFyt9w5bz0cHjYvKOWI1RSJuZLhzlpUfbLj44VMDbQvyE8VVbm1NFgZdE8vXBOfFM93d6Qza
08hFlf/Ry97h7EDPgI+HZwwBZL7ugPY0NHaQtsFR7XfxV6UAt6OFQ/77mIHSLZWkxZTzmviXtEPu
Pvyg0N/7DjIld2SoNbFvCyKtPsueaDBmXoZz7S5vq6BtMa+tDuoNL8CEN1EDFPMVko3wMubrTOPb
XZg9Zi8JK+IVOdN2NpbHo0aoSwpuYNWkZFyrQ0QziqtN5sDNZ2+duuNONcuzpWkrNaN3RQhwcZPU
6jRwDYdaf0h0YE6rUVtdnMl4XMq+kO2DV7sb9XcI1Iu0KefVg2zNii9ml7kVE1ZP/cumGobNT52Q
bIv3RGJzrU0OOrCBGg13/bTwcPmp+B9TxGkxPW5B6hYBMzVxYivj6OqNqLRrP+TNpYJKeVcIX7+g
wsos0R6BEFaxdNgsqyz+PyBnDW6ouidktjuDrZHNgszXDPg+NxgQLFQW2qwDjxEcxK+aARHkRXs1
kiUnJFs71YsLzlnDRMoIV7ZLWepJr+BlKJMuiPuqg6XO4J3kGSdSlgyZnHwQm/3XdCItwUnW/S+e
BhlEXPInq1RvsLeuLH0tM+H9SWIYJtoctjcGH95WbBXx4J8IxTdlENUpx/TjciexXZzrv3oWnJMZ
pjYh0CEMddOXOgql0QgPujJ69gsUY/h20jymUYE3vNSbzZ6akHM3TUieY3DFj8d94gYzq6cXkW5a
MoQi7o66YfB8YrPJteZ/E+ybJLVDNTT094h+zHfDZmNLjhmGgzXpzIdUbTRl9Xe/Q53py4pfJhRK
YnbMZmxYwjsz9v1hKOvyS+2jIUdargl6nMD6YT3Stn0Hi9SkhZRAb4lxjITQeKzw0Rt+B0uiPLMo
qyAyTcI6IFVwFph3M8CvJyI6eV0SY0Tci1axzYpFxxdoMmsDK+duik8gce8072aKdHfCnZeTEeSE
ugUg5JkCArwE5TXEg/mUTi21yBJkw1hQ4OdaBwDHAo/LC0fzj1SHxwMGMb691J4uxdoFBwBh63vo
4/kiGVnvo811SNyG/qZR6rmIR+cGed0w+o/Jt7MeVCLCaoNijrAeVWRVhRGcA1ZD7KlmoufYWT9P
MlS/o7Pn1yfA9pT6H22/0IZVyZAfWhnHDIcbXh6k3e1Bd3i4jf701OyJNfJXqjxt1KQXQqLf17rX
AwgGI6kMtJl6aQYLFLvKwpNcDjz22bRSepLOFaCO3HGVX/B0SbXvmYjGVAKtK2LgGlYCo57y565J
R/x1Tl8UKsUVqf0yz+9fwDuSJXb+oJZ5KjMpK8tq3mkgu/vSnXaTKb5EzrTm0+W+O2vKPpQnzNxs
8q8wOZ6MDXzp/Kt7ffL1Ws/Zp04seXn2BbgwyfW3nzdMnfwecEmTj/RnbOPDxCPjpTc7PceVGGGq
MuLvS5SGuVeVKj6b3SMPBHqWDizC/L3an67WoytTkmqdyiHgUwut0rdHsdBlO6l3oG3HmC016E2z
oXrrgerZu2P2OHA08BIsAOVHsgZBG98DOWpLCCPtweOgmiBRQgTUFQfYnKv51oO9iz6+ANLloip9
DcoIThyNnOhPMH7FeD67hV82m/dxlbOa4kHsqTDxt2PLA6bMLKmiblxHa+Mi3zH6NR8jrVg5p+yV
4gTOqA8E23VlOK7b4VIoWZqyXvvKrGDGpEMc8LNBL4XHs6dGXQcP173fCq1xfNPcXeUHbK7pDPox
6zTTPjB5o5Tw6QsKbjv1lG/he0aLY+6qtOzutSuy+GTm/5f+YgwGcAjNPptQLY3MBNZIkiBVjT+d
VqJMTosOPpOip5wmO+PoySVofqH/3L0KB+txVaKgYmnDscNfIHCuCgaG7+L0rKVyhbgtYmjsOOgj
HToojVaayFlp+4NDd4v8I0Iy+dw3Rz0R00+FD0DOY8DfOP91uHEpMwD3AoDS56B2VuJsZL7WDlYO
yyzyrwTPwHqV5IXfQiFCY7/4H4tMfNL4bbI4OnqhgMhHGZ54nWYZskG+p2oSyn74nrDZD3MqD2rN
qAtjGV6dHvSu4/wgpNwCY5uNYpqRZKgKjpCRy9gzlLYmOPSCmOIJDWfvxyPunr51/2RPpPDkvxVK
4KxNtup7CmAQatLwPHagzu4LQxkhWltLEx8gmidramTcCrrg3KS5e8936mIwv3LA4R/6fFiI2NoK
AbAa94yhiXd9eotGPLPgOJOysz2J9I1vdVDfBKtL7bSrW6PKDuTGpWpiFU9OsbxuhWGUZAfVWfEc
Gq+gEsat6+UUHirmOGSYtR91kQdtvRvN6gJwquaJZFO1Pc8xFdrU1CSaqMyYkW1ojTjGWo4u52aU
H0fegXdFNw/hjqhtLDDrsteeFVVQPIiDhKtU2xUn28WZNp3UEUtvZz58wUCSgSiZr5OD1d0cUnT4
Dtod2TtMgfEaPcVtyMH/2EulRkMxsIANmon/5n5k0mWMC0UH4S4CvoVqKQOMySZPm6lSKJXQSRre
8oRmB5Hj7KQjSN7vfiPEJ9PFGdGQjHNWSZ5Bd6kKkwkQ9En84AQv8aPSxli0XIy551rmgO55IjPK
+IPZRXtlPqeU9hhFfElKb2wsTiQr60QB3RF8pOEmfmFleYC0P3JFu3Q/dSVEA7WwAqB8VMsQy1H/
E0E9/j0yxv5ghNrCLL1NFZgF2E3O/NlSfrWS268cVptaFCnVhhkqJ5xHoLFe0eGbq79X2YEfOKxn
DA9d3y8+DrFHXPbHqBAD78nE4CHUQ09DjAu370OS5JAVG7VzoO86IHDA80oL2BnDcZMZauK8p6l4
Gig+UDkF9XDpwczGFBVXrMvO77PlHn4II5DhF2cTA55XAYDCbY6KLFZ1a6dtW47/W6xR5qquQVtB
3a/U6niGd7IBehkF9RCS+uD209fm/nMvM5SxpG7LwvaLGADh9F4kHe3yVJ8hHYb7HWoSdGEJ412b
a2qyUnzq37VA9LAH+3iGEwzia1FO3rDRSx5GfEPeC62eIjBmJmpHO2/KykhFGNvxYdc93UHgErIa
LWMXE54Cdn9kOJNa0soDXYqc0i95M/aMhyUWV5a/C68L8oMOnhRwoCIr7RL8YWuvEZF3SvYMyiGc
d2eP8ExKkioxlIs3OxnH19qXHDtzOyopbgTK44BLqYb5BuUoL27Q5EDpSisKsJLseB1Bvl5pwquF
0mBMB01ZMMzTaBWNG1gk/YfnKuoQIv/cnCcDj4+qTcrhYPBJ6dIWv14V14EjsN6j0N7rTqrVKKKF
rpUeGhcCIGzhm2veQoHRQEZpM/d+42j4AsUaWekLemKMuB8de1ahZHQ7w3gFqeGn6K7g7EITMxgc
566rKB3UlqKilMk0bU2aYyxMKywkyfvJnb2Kqd0mwWi4VbAkNoyS0h0mtKoWWyGupojx5PtiMVKv
QIEwPdxB2NpVE8jEpjOeYZAenLzXXtVHuVS67uCqHb7nrdAWce7rMpwRX3DtWGgqnLf3wM8YdFYs
1/3ZltfURqOdr3SN30tAJjRpwlFm8LcO0EJ3KdxDffEJAB8gCyjchzN5U/CaFD3TL0cQPhDjZmz8
OAoE6VsaeqpBN7JVqoW19I7ZEK/mmqQZiwV367+Zqx5IyRdfWeU6pQ/oD/ZCeQqfMWhFJUytIT9Z
VVlpMlTOnnkauQNHp1j9s/V7yRRJJPU1Sm3mjvWEgfS9CMWytggdnKU8zyfd+IUFGYoh69LTEi9F
Wf4qolJijH33b+fRDTtO75vlvCV47HnxY1E/OFfHOZpnEBCG/ftXQaylZ67E+ogfRzPiLWtweXSG
WZmMoLWCl00NgxIq8o4/jBe3E67MttGa1F1tE2N0zmtfEYtGejT52BrbKBkT8maPqmqIdOQvG6by
rClUf+r7s+Xq9BOL7vYqmwahW+ZxdRDQhlgcSOJM3sgg62SDQRmoVujHgzDAi9lRjzX8HcxunOg8
Crmi+pzaCPnD9UjB5EZhy/ChtBW0KMs7jlvqAGF0CfO05QjlwnW9ZonI7vzRX1t5QvrOYptgays0
bZjzkzbH/JDyewVryCsW3Ry4GXUNbX5KHtKhOD9q2kGlhyCbGn0X0RpcpzAZN6tgfUNtuMbMC0vN
4nzKP3UgBuYbod/neCeFN7d3uZq/unroOBB+CSUnFK1N3/XzuOfNZas4sDKQFj/4QcocBBCRA1Eh
4PYncsewuGi+tCrpiaXICq1X0Nqhi0463i85TkNKCtxsC1jY7SBN2B/MFd69xXJLqR7L0qzkUQyw
DwHUUnp2+yCnY2URrbz8BCNTFjc8YzURtwRMR2cf/46tm/d1BzstF0NdQcZDimd2aepmfRj8anXu
N1fePCrJwRRfGTbu86HTO4LSEu8+LuLI/G9tGdZ69Z0q8IvYHA1A5gLmN6A29ufnRCmIfB4ogYbJ
iVjhbwHnXn2yyuC4YxRJ4zcv8giw70+Scw2s3z6miWLVIELlN11yt9ci5+sN88U1wi2MY3R5K+VJ
MkAQZZY7eMkDj7Yjcy0j/Kx/Ku6rdsafS2c9QUvRXuXt4W36ckrbylAkwFj7KzPAN9GLxRnNz5Zl
xBo0Wg+Qt8u7sFX3tr5z+oUiNkfzxlHbb+hAzKEvQwQk0tDEFGB6XustqKx9GUvPxlHjNiGZiT6B
Z+kXzE/Eol08J7uvmtONqVpJSnpY0rwAbmBVAKfrq2QLWP9l4smcF+8b4uRDSV4YVYUUXicOTl1Q
bl7vfIXsI2mpiGdiKPlsKa1hZXIk0c2PbAGwAR+Ov1E++X03PBL7d3YEaAwz+PLwl+/sMbXNlDM7
foXyPvsRlOfG7NpzzqHzbLdiH/Y+4/rtTyIsuECKQuYvHyQp9iqUKWlTf6ki7dPlYHDK3S2kqWZI
RjP+TQIYaYy8HeThmjdWFrmMQj47u8UkNY/kn7bG8+SqLl43dYOxsAshmfBBe+Kp+ax7SZAQi6MY
fjvHt8lc+RhKI77skFYSCpCfo7o3UghzISJgDRrdVfwOcYV5kAxL75hVVdpytM/ZjCIj3vgchkOL
+9CHcTPMcFsXSqiTsQ6Dk4xBQGEdDPeQAl0miN9XGOhAPZcFRUIDAWsxT/yxHi7LWMMw3YeJorb9
0duIZHWmp+eRBGQT9u5grsThKM7bW+eWMiiz16OsRF91cGCku0S6cNUa3K8GSnMiH1mq+wJWa+/x
K2CHPnNtr+oSB2bTxdoop8Q8NCa4dxq2Fbi1qPs0ew/hE4ps22fhXxoH2UsuNO+7JxenskgYLhGY
1/FdKzhWdZyqs3acIec31I0gN/YPfpc34aXgFHN5QWTgZ1gAG4zbRUw6HjmCppl32+PhtDGZRcEP
xIsHW9Z8URLCnhWmeAiL6xLAOccDE/SXAB9y6mxZ4VF7GqESIcs8ev2vWUvJ0B4iJd94fe0lWk1Z
F7NMaOzNtkZkSIP+zwHl2XFfAq4+rQ0w1JvBIAxVY5rL/ilyjFHcIuFLXH7ef9wJ84aqXlTH7JnE
ccd+EiPU/Tw8+bE6EeTOuJ1aLSAxGkscHOhc/Wep+VxJi0NkYVxORIFWUZIiLGnB/ZW0//3gcSUw
ykfb8FS5Z/4ChyrjiTjUttVKCttNOoWfPbPcCAcFDkoNYVAgEahFGq+dR2Fd6iU0be7jaBYWZtOX
Xpec7zk71ga5U6f2cTcMl855YFSHe7KgoIKgXUwYwqzGw7/aTOTe4jH4bXOWdiFWUOvPnmM7EHbm
NdjWgV22xca4haP/Pzz+r3WoTarjQu5gtC9yp8UjHidMoNGUqvIYrbVOzm0N+30B6SaITvC5bFeI
SjielmwML/KtWb+4jh7LhVXEyuHORZwVFPnBYIg/arXgS2UY2ywbBr5fSc0iCWlAZXFf9xVz7eid
SfAEsTEtBXvGk68rDCCmf36oyuDbhQ74bB/NLeTUzNcLY0VSmdgev81+kuQ91g/OcdDkEgSdA/Vm
dWpM7i7vIbeK4sJ5dKPA/AH9g5mQ3RBuGbre76VNm9wAC9smXx4RUqfqIIqqcOJ/mel948kSIWAP
3JOKLapdUcoMQaZeb0akdgTdy7VEAeZdkqO26kbRZcl2oKNcSYKY2YBD2S1jZO/aSvOzEyYm8LBl
LPIbbjul7z7na2MhnHdEOYPN2ni+D2F1MadCyIkJtSiLrdKshtddFRmuJ1ZU8+RdL63kEm6oTOoq
dOIJZN+lXIz+C34shg+KkFy9NWUP0oP14Y0n4ehpZx4VmHbxvQIdYQbTBmdDETh1uOTuy2YMhTQ6
qTyAlUwmpiBqfFWTU2zRAOyOO6wp8ndhuc7r72ehKa+Lwa8w+qdaNkVQIjjAJ/korVxWsvgKMzhj
17ix962PjIs8T7Ao8P5m6LvoFjNyHNcOLD55Kcq8FPSXCVJ4HnR9YJOd3D722kKsnCCfLb3TfyAB
3NNrVR4bHfgaM+A+HUwzgU44PZYY235TmR0r0/RYuSVVYuadspYmfgNOJg9M2xJ1pACPk62mBevl
65yTpBHcR19+BHV2r81AxwK3MA0iTNed7I530WdRsC1ks9fhITX6WyXVcQy1f86sT14kwur58cdC
U4bEc2jxBwBNfEQiSH4dKC7FtaSIXTCcdgv3aMafseanU4LGE9uTIBLW/DwsQcvZhC+18d62MUrV
FdSkzRPdzQtjw2KFkHcDfSEEbjhu0bU/Aq4zFzsNkUmXxfCXG1zyd6Esfu3mHyLbXPzEM8f0b/F7
vv9Gp6bEPnm8OME2jy1/oh6QDfRH5Mw+cXAPBzqo9m9wnh3ExY8AFMzXpxwruGjSdF+BqFZo+YcM
CgsPFTOZhXdHAwc6kX2muSZ2LMbkFZJck0MoQeMzmJMpn3JFw/5KoDdA/GHIPo/n1YyNDpibjQEJ
ekuvOi49C5ktVSPrP0QZpEsLNECSpc8uRC7RRDnoUbL45ReBkapXw41fywOzmjgkIkPIoq3wd8kW
mrsA8FcCcQqpxue5fuyZlXOGFbN3/glFBnE8qFxZJ3+VV63UbIIrosgQNS7uXcZreGduALuggrCt
3PylovapV1/h+WrhrKGgvjGROFdbthKR3XEkUTpvF2VseIMfr9CzBzgiE3c35gdP0uurGmc9SGwe
iklGfS0F+ByulSIcJFaA0JvWE7C0Xy1XnL355wb+ZTrxOex7t9LDChnxxWlz0MKaDpAvPRdqdauV
RzW+zT9MzIK0ahktNpifcghjTHAPOQvelXWS2SA4ljOar0uR6cQRIEHpLAdoVdX7V1eyMDH4PZi0
Bv0PhlVSRl6cx2suQzOvHZFmVz6GCpQ3iFHjGzmOcv+K2xbCE5GOmYVCTptGc7Ktf94HNARnyWi4
ioJiC3kflMumoRjPFKpcwYv3DtRecJ4pcCj+n8Y7Z5O1pBoP8FPuyDgFjZmTtPrhWSmJAUB65eXG
bDY9zlD7PDqliYywXfUbivecfN1Ouanrqb61EAqVJ4uwJc0KxIKtYRrQLN23lcJB8vpDB9VDss5x
X+2w9uzsHWfhAGwdz4ieIBxkrr2UrfUl4A8pe5uKeidAHtuLEMcec1BV9H+YBsBiIF5RvRUmM6iQ
3qeueJA/YkthFVXGRNnCHNg06Xyw9YBPlgFsA7Sgr3gWxWnyMol2cP4LMz0IyeB067oQlht0ZYX+
9YO37gJOHU9RygGcAUZ2caOxEFyWPYE7MHBlWqatggQbs35nr+c1YUJCwlllxnfV2G7D/P6AT4zk
kWtKdyPjIsumv1Z9KUIrTmN7qWQx2mTyaoPk/dOKE/hCogdcvE2qqPPw/FIToMHf+dVBlJbfaJcL
72f1C5Cu2+nsr76Lt7cnnCRYaJSpTc1CW2uKXhbHEf97kfE0JTDJWPOW0HXKVbV68odNElbTVYQz
sbndtabIqJJ8StPgXzkC2yF948dlVdr03aDXMvNkGC115P4BMnlvTKvKu/P15/Fq+sV1bnRrpr70
Abm01YHtJSWdRs00+r08G/D3bFNBXQSKZ4MsuoS95aRqX/ItGHCfEDfL2BZiYusIFlksBPEJih9o
DTiJaZ0PcCUheJbmXUMt6C+YsHGIntLhZ4nQywds5GC9Ch3yWWoB6EukjjruSc3uzILlNO6yN+n0
UfNRpqB+myJjVvXwzeltsq5+bfTTGVaUQWqCQYWlvsKu+jU2MilThV4+O/MaBtEbitwc++M/10pM
nNYTs1Q6Rt3m4/7Fz1i15+Fa4D7cdK0y9vC/7eAJl8RlA+EAcoR9z3IOElOUKBC+LC9LjS0LFI87
urewlYwRtsU7IxGDP3UYG+/n2+qPYUzCVesWBRSkmjmYOPbQ2u7bl2VxgAL/e4D0hUfFhMsROBZY
/FOxIqUerqJVLIu6+QE57t7gSzSkQUq85xylum5FK11qrnT/vxMfPbg4nnXv0CxfjeLGOIppzWWT
c6X2QphhYfOXSOeeNslNXhMfBHfhRwtm+tgYG1t8PIGIVN+lL2NR+KynM9cEVS4/IF0UbFO3c32E
iEKu5FjDdR8DDlRcqYOtkH8Bz6ABifLDV2FoI4FzLfDvS45jARaDA2YAV1b6uJ2kwW2fmdmRASpp
D/RJ40G6Zrou4UJTB9DuMGWCZRyy54UpsYcfEK3LH9d1wXpvKv9L89rAgtqR3U/DWMSHYsYplgHc
CQNB4Ef7cOOluh6Y5sIWXraujTi1O6EA3v9hYkS4YtSCRp2K5nf3PLHTaIB++yrHtPxKkLYRLVfo
xUElmYcHFN1jMVEs83kwlitQuZmLIsRO2/LVu0GG0YZT7oGhRAigcbtcmroMnWZmgcVFoO+o24fW
t+BEB1/mbGtBKu4Xuc6owYtjBzUy/8OVJLGJymB2mR4FChlSlErnNosGtXVaLn6hK+7a8VNIypbH
EYp+drzz9WECZt3ttbwBaqUku8J2LpreX8Six3WnORHy50RetAXNM7I+mvdu2ZLs8binquBDa+Q5
xZDOUpJ5rah4KRO1s8H+lQcBNPxajo1aqMaYGOZbRuP3KDjUtk5nTXfQ6WyhorBTtv1AcjheJMGU
mdwvqVNvm+5kSjdEEN5ubHQ4pGns4L7/vYfxIlyZ/K6vOPaJoL8nRIucOapVtZ07SObOBkY7LQQA
QJiVHxCMO7/atg2Pvw+0FElFkkJ3MRbGO4feEXXtXqK6/0ADvQxlviRuLQa7OmgFNizGYQVTBb8n
FKqZdzzHuSiX1AMwHNLrCmOZP9Mq3Gq5A0g+ckgt23yoD1VmEUFiSZslayBxLzbaA9LGaXgik5uC
af8dHB8d/lqsfOEPiuKlySdDx5f/ZCS+a9VnDCq4aTsPjE1zIo5uE52xEbJobqLGPSCkO3BOZlaX
hWsCRaaJkILbD6pSzpqUBQUcfWVqzp0afsS3jtO5siRu8iKdDWzD5OeAZtiedJws1WMxhgFQNpRs
3qNDc8NYVUmpUGjR47UYkdDvZ8CxKrLZRh0sP+FPCIMmWT7PArQ1UC7UeafxrV4rGVBvJbLXPuXB
Gir0vIi2KJoO2zqEPEP94vKqwinYweO+I+lOc37WvHlvQ0piblkhHBURBxqB8F0VMUQGIfNx72I6
QytWhLc0LdVYylIo+pcBvxeXXDP6ZYnDphgfFKcPtrgXFSj49Pr5xY3yuAdubQPYdgK3+ObZ46l2
azi+pRhrnnjsuVZsVcLfWmxqY/ruZKUb1mlUzOeH9sGYbCyZ/NROt6A2Qxe6fzSFNcVT3hJ7f0uG
oXMZofe9NLKuejGK/6kYQaAdY5sTRq69WG5LvmCIa7AnIQJXCdqPzWJ+wR7Bgn2kC664xkd3EoQ9
ZSCCFcqgjpbV1JloH4Bc+ihgrD3+l5L2nPjgasZM6zMAVDu2kedA6I8Nf5RGQuZ9gF1zUPiC6pZ/
fa8zIRb4P4a0k/xgi3RJS2yLOZQWRMfkBSIy/1pUVRXrrojD67yBcoFRu3Bm8p4Y9Jn5hR0te8Lo
LBq+COWXnuMBQQ3F8qNYxHkwN0gDBySmpYpKiW/2JpiZOtAWUW/n3xd63aVIe6A0vIngfIhZIIMX
QdUQw/T0Ze9Zm90gKq7kbaAM+ZLfnZtq8Re4USrcGH3L8/IQ8YXXBzIkuq7KRAb/KPJPUXiR3x5R
QsOXNrGKazW9TLBipJGfYisyuMZi9VUR0toDoDQrDusPKQJLgGjFP/HR/IRoR/mdbdUyC6Vr0GMI
F4BqtFK0AT+3cxTXIjE0IqTtbyIcRf8jSzSUwfL0eYv5L8iOnNMaWYlj6vvZgdcqOxM/VFbNcZT1
IqgAbI9jSgRHJn3EXCJsUvpnuba81kGyRjpcgeoEzOpbUZSvpyQOKcouX70RxiRM4B/i3m7feNjS
oa/VmVvr3yN8VQuefdzpHNNPrZkiX0YJ9z+kbS5gD6cMpEP0OPH0C2+AHE/BCp/duC1jd1SxMydt
50WsC06bl9ZH3PVUvDMGOy5HcgkhE44S47BatWwVvVUzgt84Ch1gqcYw8uhTmGQzeDb6WcuGcc3C
nlydpD8BaWuWALxlW5Rv3b9MobuUaluB8yP7hNivnLOK89vPHjTLwp2QwiWBZL5M837R4+EYs4Z7
A50UupBAlYTnKm8YlJgcESPhb4MA7Y/n5kZX6P+eoUoI41NHjLUULIXVwE+0SS+CCr5mjZavKd3W
0rTBq5QAdWr67s2e+XVh5Z9fjwOkjVxaRuO3pxSqiXqo4dhH3qbhcuAad6tMXNyOW5OTV2euWvx3
nMoUtYLwLsmA0kFIsmIACGYLyOI41oLAsetsFmMMn9W6jw8SuReuuOukeChSgfXCG2sSMJCamT2G
sxoVbr4O7Pz1w/gz07oRf7acSTzwGxeVOEpzJzgzMRwOb1Yc5NTEJumzKM0XTqaq96BnhlyEcuHt
43Hq8UHV2ntdYeGy2SUI0aMdTj1ia4c0vtZ5Bq2tEX7UZnda33dq2U2p3s7mMzGxG5Q3/iYXi52/
KlFfU/X/1f3aObCu5V/J4+CosHxAh3O3h7fOT0d4PlWeatwXsfV17r/l/EYnGE8yLsI82CDAFuRX
v/FgWSjR4yEQt776XPh9WWpLq4gSU1n2O2vOA3L9EMAEFBQNiyb/0opA60wMZGITLc0dWoJJwHD6
l7WMjg/ckAqRWJZu6OrJnnOtezYoW+lnxbEqnbLLZMf36zstLDguuZSThPSYfqw/osMubzIePRGM
eV1fePcweDlnJmqCaexZMjRBuHIDuGa6UPwvyHCxRo/w075bvq1NwSM4aYf4hvEW6mgq75qeboAl
MTBGiNnuzpFMsPzIGLbPMBU2CS1Wa6vXa9yb4zplTsp0xVp4ajHCM2fm97BsC6ehgL1XsF4DIjs5
aWnyU62QXUkvbHaZ74xceOzhHUj+wfpquGlH8prj14UfhX2ImbyVTCamK8W7u2/mYdroGaFx2Lrc
wSHrRzXBy2Yp4yYigGIo189tAEhPRYqHEx2ys1K3q/yzlL9RdcilRawKXr744mRozsZkQL/GH2+G
8ZVuHoc5Sk0lZKoCbZ8kxgqChguIz9NSRjDl6xrLnOJp7bjxqc7n3AzLtmZqBfWxNaqxfyMqwKae
hDrWD32DHESmVS/naUJR0LfAe0KzDJHYdZ9oELL52E74/0jNFS06z/4P8r+//YrkzEO7Iht3s2Hc
+tyAbzigdx+jd3ORDm5fPyd9x62K4WYecaDHp7Zp0bxT+sjPK2vPcWBvZoMNCO5V03Cpij3hPB80
SJphHgkcgRnenTdJQdI2xskM34oCgcrzAo2g+9dzzk0OnKbRGymVqdMfqke4bWl3kZo4YMmez2CT
QzUoFxHd06FCqygoQ/S4yTN2ykdDGiqIqlwnQ4rwRKq4oN5dcPl4+55dh7sTa41UoCIyNi8SzCJU
d3JQS/0p+8vj8zi+17GLLyD6XU3ayl9pZCb+AZcfKwZT4lJycmiwQvr2MWeLJmAEXxK/Yvb6WJQR
mlBU+SEB03y51qgdsDpGqmPYuG2GGNwKhNtkM487EegV1WcLZ0wd1HAoFKNubLqn8ixH4yjQy4yw
igZO/djWv80VrfNVYgH7PpLY6U37iQnKRvid5zYTBmyh+0fiPLIuZn0K3DhtpzJefMANfbWwkSNn
GJkj5uRFFh665aayAQIdxOkOvYisRomSwQjx07yRO7wG627ClKofjbKWRf9A/Qx1B2zLVn1XRlxd
0IFtmAc7Ye2I9ka+Xcq0GJKJWcOszDszBzKbFgvNQiQ3si4wDXQeSarORXWilvU9FdYy8Dm4X9zd
1UC/+N6O4YcjPsJ5tHFnWliIbpDHopesyPo44hSZ5d9FzpkIeVdatOXBdAZ2JKZ4B+jMpX7ItVaE
yLzWCysLsqWBokUommK5BtS0XCBZucDx4aLoqHg1sIlXgsY1R71JqEa25D76FDz90xHVNgUBCHNn
ZSWA2TPcPckOYnTwYOL1dqIKVUZetjG8GlyWCb57RLPL5SjH1OxrH7oXz0N8qsDB9pMe1qEqlrAR
XjEuq1betWCnb1zVwcky0f5+ygCzbl4TBFfcb2YknqXJW/JMVOkmg/IYCc35BTRWBMH0jAq73vAr
qA6MNILVLVp5/h2oDP3Rpgazue6bb7ssNhm8q77tNkxL01j9lpavwBWm53l16tK74YVev53eTWPR
6HybiQZ0i8TRQdwg/G7eNdw5v427oBQW3kE7lHQhjke1At4nKOZ9tGH2fkjtNm+rYU2L+GztGYMd
Fgsvm9v9lAWIYOnU1OdXckb61ftOmSUTw0WJ4A/hGvSa77bQEQ3tX6ZVEg+iXR8e1GZhA7JsKlKv
4cNF7QK5z2XhN6C4659tTQCPdJ73HG2cmeq20RzrZpVR9J9gX+GJSomUuEnon7ZixjdCMGRJz91l
xu6cP24q+t3T3C8snJ1NboUqtXP76nqVxBR8jMDhAdxw7zjbYO+bpR0Tb1GvbkJCiz8C3v6YQkcq
WKCU7wvZFWqKkFZ0ttJzRibKmiueaTXyahiqen5C3Ad6ArZWyqGNPg9W/SsEyFcoVl0LGhplVoNU
bwn5wuJVLsx81sfzjQ8IqTDeJySz4vn3feTDjToe+lt5/jyUkozd3u1izwfYMiiwgEmzN73Mx0AB
C6OcZIwIQTeyViLKxp4z7WORz1X15WkDxBwvcxGgR6Mb8LT3MycXK67T3EPyzl7eN4lq/VLe+cas
JA05KC+QOqQAYP2yy2u0u/nz7YL8CNgbXSn1O8p6AMd8msjrqF6TPgEAxoYrOb6F7z/o2wQCxq4K
Pr/C5oU6FN/RdT2uMarokhDnedwVqbvLvi4pMRr3LjK5e+6LDPkomTPOSjwLT44v72GKLVC2GR7B
pcEspUpvjY8fNPMlJBMIlSAIRmsiDFoV1s191APj6Qu+rJqJTipbuvUUxaMGNbECNGioftUEWpBq
RSruyrpkel0RU/O3pnnTmHbpAcgJ/LNbksOFNJlCvMM6M2TJWWbx1pCq+ajRyLC+VFpvdhw1ISwT
Dy8EI4ea+XwGBYgUXILUdg/zvmlLzLZxaudzpA9yIza1hnnfNK4Q5SGGFlsivi9nd3R7InH9UQm9
9YtUl/VWYqPyv4Y1MfxBiF7pqG/PNIAScC6INCC7AOlA7oMzCCTzvNF9zYvnpZ6CBuFyodikHR7F
SlL1ENmbcSS8u2qeU8NEvoULkDJWXd+FwF8LfBfxTBuvM1JLRMVz1BfTZItmuaPxGSPUtCzIgZW3
fi1kk4TC/DDcKRBpj5oMZ96SVWdsMXVojG6j5rTk/9SJQiKjboBAwmUNn2MZ3OdKZRbsYZUQiPwP
P/UV7fqsVPl69CDs/4ieJFlk/4MHFFZlynrZHwnKLuqwS3FTA1sK5BwoUuzIN5oz2CVOOElmLk5I
zdv/+S98hnLgH5cQV4k2i/qRLSdqAM786P0zPPPDA1cSHNDl9Z8eGOxl1iHnb335NtHsd1WrtL5o
SwbXoPmaRe9M1gdCvzR/MqSNIEuzbSbIXZb/0vxIHl8oZjEBJYLG0C8vDvzmXncAMa3cVz3rXpGt
R23NprvaCM6uehGr6zhkQELCFqZDeh+tuLcuNV9sEWdcw6bvr2tBYCOJVsdTxOg0allaIqmWBgPG
BQUDis3He3XRhY9tkV58gWz4KLLlLW5NNyl5/AO8Q+iN0G7A6OeaVpqcX+UV3o6ER/EAouDsEydK
M1DDFq8vVGp9sSMJfX1d3trF4RFJkCD6cEQMT9/eahqm4PP+j2tMY31gGqXk4YjIrD4hZ0PVpCtf
wUQtBnJd2PMOVrBEm67qibLwyI3Nm3S5mFtZlw5LMPjwn4mGShkGA/WBPUf/O+pqrfFWpN7+6Qj5
Vpju6Lc0pWngb7hH9uiNWwsGszvmBgcIoaKejVkj0IVLMVdiyWFcFA464av4tdUweWEI7ze7XPOl
BE/AQr0LgWaPDguo+v/xHXiuFgAqVYIJkcOHIGj68kcPNQLeA7CJrzqSc//47kFeMBiqC5aTUuo9
KwHDE6zz/ODHwdZYJ+01RVwB9DchuM9ZY/uFYFr8Iw9Ly4d8NqB9eSouK0wwWVN7Ag9Zjs4hR1/G
qQwKZDqVuFL+c4YTrHVGUTj9EfDXufX7qTqK5X+6/aiR9h4mAKBqOoeTHpzR18gLY+b31Me55xDV
cd7aGE5M+0tianBOE81CtDaoLeBsB3zhOZzhjAdDjom0ncY3lT38jAlvUxhRRwJcd7ZXPY8Ho+jg
30kGKIcbEZIg4kM4nAF/dNGGj7nWRr6/UZZlH396mvw3cut+yEij6yBLJ6K+6cpvnS3Po8i7y4Pb
irfIOSoNUMNj6mG0txr1eibzlMK4uZ0kaPUwWuOg63PdmyAIiskXkSwNvZedxEKi2dx8k5vAaN17
cSTzmC6EXW9pICK+ee2R+ovmKSXWbIITW0tZzQ+jc1yqyxTn6Zpl83+NYOaD1LPtyWPIr5EeuOb8
2+5NFqBuUD5YzLIwugz5xXfXMmhhmQGYm+ZHIEc1wlsson5LwkdK24SuwJuPIz6RAnLdEdxa/e1E
yHlgIYoh/3IYo6QOFAAwA/JPpg4m6/03vvT/c9qdhG7/c1/hgRaBbxsjqfJJZSwZx27hAUYK8rN6
ptYeQEDjN9pbmlTPr9y2wZtKm+9VMeywLi2xdOJSu60e+Na3EkGvcGIXfNI4ZICLCr+43bPNH2mT
EufKrnpiWZCsIqcDtYN9SgJmyI+6EfUgHRBomYnqZFdUVXhZiTQqk9Fjz4SGnL7j92y2f69C7CfH
dkzvlV2KCW8Fxtowa8xVhCuW2qvXnyC095eDxwW0+BBl2tK9TjXgZ8aSfvtNuqbESPTzHPTHMy+1
SNxCdIvSDhe9rnco9TB1S9B46qA1bpDoFaGQS/jKaPAi36wGz9BqR6pBilIkjAIYuCk4X+FhHIbr
/t0zxycT1+VlChled54Dg7rIOYZzMCCxLdxAv8Ss5hDSnS0gwPcWaZKYz5a+GUJZZZY04m5N/VHH
gSjHijj7spy5LolsNybHtkARfW1wWFxkgeDIBmUkSJrOzOXl5gDNgd7FAcXcKaxxL5iJFCIoZIP7
u11d5iFk8PUYyvyg1CxtXGtOO9rfnNQZpRUwXbpyVHttSCaOz2hWrDb6nV2b8qP3KRG+PKKJQEwR
msxRpvmxszntP3JNmMUDm7mM5qcR5zcpl+hwP2ffD4f6tLx9VZFR7LfpjVzrPtbyA4c0Yd4m1P5C
AXve+n5FtNuT1LHcQ8zYaP6vZUURgz6HndwcOJ94EHrArJ/48fKTsc2EP784XMqyV/PNHV7uiBxs
TOcBSTHWso65FZB6SoIP/3HWfQMx+/miekvhMaINgjK/3B9danUqOhxUMGqQh8vIdR+neqnJK4/3
eDt/C/tEqt25qexS4CMr7TGNP6lSgOKiq68oVNnn/O9/PUM+06Xmh7j346SvQXyQ/U7u2g2x2TPw
BBgvRkiXnNRV9X56vF1WpGDw2kXbSVOOvohtJVHGK9N3t7zb5NWDV+SEZn86TXbRaguZwEd0ixO+
JFmqiErlSAuCBd9kXsn2qpwafHM5l5+fDFfyQuqHWSX81Q8s6aeL666YwRGa7Pn8h4WY2tqh9m98
d614D9jUegtBM+3dfk7LbY0tTzBU/58MYVO/7Z+Hap2VBVTPwi5hY0yYys3pyq3JkStiD8R5qxBX
35SVgNIei8nqOztTiu/ANLCZZGRwl1PagR8Ko9X89ZYRx1uw3lQE0ul35rmZLaKjc+RNN4bjeSLW
06AlC7Qd57c3e+dBzu/Qc3LJrkQ7+49gkfVljUnH3DVfu2eFmKsmjLTy6iixRzaXVc219NE8BoXY
/VEVpfhkdBJ5pSvjrl4Xy0tpUb2TJnBqgXMgNFE+sW5WGnYlLY7Jl11cq6tEbMbqnxQ/kavxTeHR
cDCxn+0UnUN8dpi/D1P4w8CAMYos3kDO+ineZwuqaVFXhd9FNbh/xYqEar5+SxESLzBQ/njIsesZ
Q2DEhD2Rbr0TNv3SpN6JF3/YI05pnr8CE4uQ8ZDqBfcAlFY77Td2sKLeHYDQgvVWfi+Kb7GSXiOM
JNkIzIBlAQdyD2pU0c2rvKutOQuf1itF7D1RNq2DKc9hJHd5ZhMJ32m4qsCKS++bCheNCph2aY2C
fBM/EuEtXJv6H+xA54VaEpN+iX3WHI3MoW8nnSCeoX5o0D5SYbSTzGwJT6oe2x6pSveyfYBuvewz
GL0bODzwaV5P3rzZjxG+t77faTVbv8BbqdEI5FoOsFMKK0e6H/ba1tJzQTH5P6KqCySPhNA9/5E3
mAkB3MfJksvgjnxxyCqYk78ZZ+2CyLV4H4WaNx5Bnn/5GWi90EpjBzvnIKtQ3XTMIFF8oOAG2Skl
AVzuwdWhgmAQCBbEw2tJ+eW+fePP8Iyw/ngPjbCv2hl1Xu9YzYX9d4IXFknTUWTyLnZqZKgEHzKu
e7zbdC2hoJ68/zIUGVGSeXbSvkEKplwV0gJ5QSBJVBs9D1hilpJIuDi0zk52IzSJj74q4ZfZUciv
ttIwlLLpnoWPPnLiMggeJKA4YcQq4dz6RyTuYknBDTKWGxXvhe5LmIdxM/LqxuSDs+QgvU9Swfr6
92bFSr3ldPHE6JHnKVsIQ9/4+dWNBEgbU09aqDA/ejyBhoXzZTFquZrbHmbGpCNHhV4K5z3Dw1gL
tA0PtdLsvuV0Ki4oYvabP5JdJ23gQNlptuiJlSy3qGSnt37eXKnMkdXXWOLlNc7MBKrr+n5nyKN8
BOvgW8w+NtZ4nO1INDGr4RAXSr5Iz5QjvIL+xGnsXh/nrFoOyNg2L6l90n6FTIFN5QfKA9mVaynd
5oVkw3TrZ7ax6SSofu7Lubdf0p/YOOHYai0b9DYrb1xW64edi2RrxkiCqvmYAE+5a5dXsUUYXDL+
VhQa5VVpOdmU3LnScfwNTQm7VGa48i6k7H6LuEKSTJ6wfDEQqU1e0j+lSL9XVHQDaUEp5siAIimK
Fu+7OS799X/Z8gIy8qM79/t6qPcKyF6NDBsMJ+mlU+uI3osdAb38lShe488+SG54DxUumD+7Edbp
HE8AUWuvjdsWo1cXE4+PeIh5GgFGI3mPowPYD/iWSZOo5wdKmbSYb3ehOpEArHK9rLbe/dpc0FDz
p0gB5sF00y3ji49n1kj161X8feLvwS72iK6aeX2n/p/QEx2lCiVzHL5rUpU+NQ5iUymPETv9A/An
EcOq+N7Zm5Foa/zrFQJDQfe0l8iukrwNYNEevQxGSVyTFnPRttwR6V4QZ4ljbU9YiyAkf64GYYIM
Lp+Bg3s32FgK6JwRXlQpkMh8D2/cM20sAhWcqJJbBfv4wNsf6FvpA/T7Jvnhb78wExmtc7tf3DfT
f0Id7GppbsesW5zDrai45TLisrsMfPtVNIu+rKoBdqiBSsaku9RL2Njv4biaR4HWEudF5BgEluTu
Ogv6BNqp4Lrx8RSzT/XlJIq7RHM6Qwo/G8HDcqITOzGN8E7DT2wikuJdQmjWF0o5UqLgXocwjylO
wUSI4JWKRXb0tCdIhE9EgtlXmjAv/DXfgBngiMnVsMFy9RH0EwD9izDx0cQi99iDyp8UF76mSjMa
+1EeGDhe+b8serg/HNWqbiYth6gHlJfuz4EaIbbtpf12Bfvug3DgbRo8xEiV8rvdB4upGOl/4rzo
YvE1FRJYq3PvUN854G3OrEqgS1CzPKR67VHZHgLvazbI0y73hv0eThAXxv9enPEd/qC4w6kIZjrH
qfsuhx/599XAUmWzL60Zt8d8w/YlNXKNH323mrZL31C6XhBZS+gvzsjzlRXt61EbtTxbSi+S+c2O
NZDy/AMrCzYWWGitzqUTOHVmrEYqOVEdRFDWf0juYF2JzE8XXFpzxJLVgc6+n/q/TjtqS7PXOqg/
uvN6sglCpkyly+9ib4iwDzlK5871ak+x7UVKWdy8wKLsWd497RXkDvpXoK6Q/gC5rBwN97jCeOG1
YtqMLOSSbOhVKMt00W3othOmh+EP0LbmZZUVQH4Ot7aF0v7qRVxenVImEHRQ5REuuJ0jVR69/p60
iYoPUFEt6xTnJObHMEAfeb1coUl7NoL9RwO8YwxoN+h3+22yCZFldBKEuAXqy6iuPDy5CSsrbHMg
8TaPFkv2nsRmYX4D2VKmLb7ZD3CSH05Qdaltw+tMmbuXn7N1YE3HHKCkLZua7xN6KkGPsntyDNlm
fsJ8OL0qBYvfBtWOEpiJTxJGMZeIN3MIkneKPje5AjYieTAtF1ZuQF2eYjEaIHuBFyS3rHeQJWiW
k3gIkM8nVmeNNiNyKVxC26bJmNP7WQH7PqalQnD5bo0PojA51qewsaq252SbcjBCO0Zf75JcrxBq
COpqE5NwCUhOuVrJqqFoTVeNfxyMvDlD86yQUXtcGWv3K6VpoOQZynUNs5Dz4UE5Q5VKIQDymMAw
mIdnkbfplPu5X3rjCO2pAmV89ESFnnuf6p2Savq/b+Lg+MKK51GupY1Ldadgv71HvctUHIAFL/Yd
vNh8RPxlAX9d2hnoy55gl6Vdhu7/9UDRwp2q+cqHz8SnDq8g7YXgajxoJhPi/98v7bjHpxdg44D9
Cu9O8kHda4wIecHp7nTcj2PTC0+7ba1lqaeulj6PHW7uncl0Tawn6jmR/Xj893V72IjOZ2o1Jtmp
YY3kXIuqUIGj8tbLzt+kl5ozK2QFCwowiYMaAZRXNdVNwjo5MhgZIlLWcT/0oT72NqkUIV3butYZ
UH2Yx8njs5hjEHGykSLdK3Hx1L+l73q1hvIYSLKBCyTKUkoY4QI895QJYhSRn6pPu6lt2jQRcEV1
CYuYInjyHfiY6CvBIxovdkNIyOp/myskY0oE0cgaYbjs/UA2RWuZzwq9pc3sfXo41/WPgOHOJGxc
TDujZ3JEev0T6VSmX/PJAUgugj7HPjPQf9lrZEqmgKqtIjDB6RZsTxdJ9BC6BZ4s6S0wb73i+HY/
LJtPsPtvTfXnpEZXbka7Qsqe2OtDDZPfByAbOn/0mAPlZ0eJqNo8ffGCR5yd9riLfpsYl9+acEM1
M99uSHVnDnk9avQsGsUklxyUbeEOJ/JCDFlOvqboHu9pf1gFadkDxQ3B6pv6fmJfbwo0Ub4HZ+Gv
x30atsY7cYBfjUDagZbj958c/q/ASPyqqq3f1L/nfIj3eY7lSDKsRc3VFOEDVbBDX5KOfE9uktoz
txyo5lHGdZtuP8lUZ+wtlmwsZi1EQKwLEHIpO5LQ7+57oCfvJFTazDFzPoirLLtK1YsYavwXVZMF
yIsgXC9tgvKot+qYtLrg0c0ZBdNm/PlIEwZJL21XUpp3YGe+yn7oQ+3CQlTst8fyOXDKCnAsfsWt
9NuAPcHDlFk/c7U2okSb1aUUNOn/GipcVMAGNct7o0jBRI5mZHQ7GnN7Ul7m+0fVtPP4wvYGw9ur
NtaUL8iBodJGMTAEmRyEeyJ0GnFkra0thKb5uafdpW/kUD3DGDMsOnpN/KEASiqJu96zMeqyI4Q8
f4y+OKu912t+Kv74rdl7K4WgsXHA5pNKdFQiZMQr+4cN+hzWEQKIPvnpafzWMi4GS1vZ1HndVzqH
8bPREc3ervRv9LfQ3df4lFxs8idnyMIdgMMJzS38/XoWWyuVymzcH0ehr/Zn3OdacTQN2Zi+Jvwt
2PoxgnXRmk6MW5kEVlh6BQNSad4NwofTtGgJLl0WTd6C16oduC+YWdYbfDLXQLdRhhjCEanYhN77
hVYBkcOhHSOrel7a/M0rPEXXqHcmFjExvyNxtQ2ka/pcJcqPFJKHBXTba8VMvaAtawimFoP4SeGy
Yw7babR0w5jvvypTnrd0yStZ1+mzKrctzYQlQslOPPz4DXbqeQq0KARvkExtBchrimqZ0u2QHxue
hZOvkP7ODKu+bXJFaXKTPvphEGHKttfZk3jQOWXT+9T9f0CBoYx9evSg+zMVA2HbDajwTUbM1eRu
VDK4Oc4M/Jom2Fb5YiW8YQ+aFeldTTRSsgvAEBDiGGV6w6QF+8yODm5Rvqef6L70W1TqlqOClxVx
VFkxNdsSynLggZpYQcTZDCAdmPQ0J6/h8VAFbusTudRgP9ylCs7UCh6HaYK7I8Oti6Zr/ccqZFgS
Of2dSzaSnvq0H/z+PwNrVlNI8xb+7osUaXgtr9MbfLKKsuRUQaLoCiOVTT6mZaK0V7yxuaH19Zoc
hcjW817On2Hppiz5dWW0kpkCjRd3KSvCelyuI+xPP4k60W8KdoPRnRhIdWjDVHvwHUQnf3BPjKfw
yVynwrFIe8RXyu3c0LT/vWI8o++qe5ReeVhiVtN/Wxx0GoV4Tz4/n/1PtUC5NV5aJrrjBRwtdn7a
Qo6RaW+bKJx2cmRRpu99+WyKuFcayt3uWHvNtAejO3llkV/0ieNnrTOYgEj12bFWUI7RUbZ2tJH9
1CzIFu4i8Yc4vVTMCtMZbL8urfV4VF8SWxaIc2pbd+lrKTt4YkAthYz239Z22uNCc3ABVSTYj/a8
sZxaaxDDUltHiFUKqsL4KH3WMcgfiHe6Wj405oFdeqdg2/b1mnSQFqanz4jNEEhaBRrBC4SZpObH
V3XqsZIr9W56WzptQJNoQUTyo3VNgbiQF0xp/OzPe6Vrz9tDFiD2l64etuIrKFHML4uA1xbOi3C+
JJGwhw8XExpwf+WRJWYJIlv/OKX3WmQdnxK7egtI7uwhsRgno6R7KNNs162wPEDVT/rzGuybSu8r
1XVnkmxLZN8Bd5c9PmMZ/rCbyfn3u3CAQjZt5w4T9/22uzMIesNMJ1N16SKcxGRsZxbLK00XnqzC
PXyyf2L8HKo1pRNmN0UstQw2Y140Clo+ILDJ+28HNWNdxGXkTVhadLPTn8S8oaiipRdbAPVxhcqY
z/Pxwen75o3Uzu5Ng1tOiETXxYjUNQ7ucLYnce/3F6L6S7wdp2R0BAjCDxDE71xq0EFaWe5XYWn9
JjmfnT8YX/K0IT6qizlxG2p61tJ4QMlDE9QRBi0G+a9EHcbkMpduS5YSuiUVfWWsTnO88gKP21+A
OHL6Ue9ikUUyimqxItgxWwL/+KgJiSat7A21N2/lipn7f5wXhsk9LAsu0RiSXhkaYzsLEQQJBwhw
zMmDkmzl23JJJ4BPWqcH5sJlWNy2ui353nTclE+dk28wHiA/EOx/57G7A1W9DOGFpJX7ignmd5sz
flmNFyN7pFhdyMo6gnjniLmZB4A9ItaH6qDTtHOjw/kFR1wgnTW0BR27RRFIEju7yQgwTba8E/sH
VUyrMSbVNDUkdAaJ35X6SoWkWaP+0owySU0Ct//8ZDPE0QaeGvIPaP+psQhoHlO3SQAyUPedIn/U
3TIJYIrqzUB7w0BhUwZwSbVou4NW78/DuziyeOOdvG/6xVfaIier+4lz/ZetncRK7BGJTlwJKeuC
AghnaksKgoqlBwyJ0vzq5gSpGwamLehWPSCxQMHzO44gnDRHTK1/uA/tcXs5hpkQQOZqtuZfFZQF
fIMYc5GwynBUKsLMoZ22EFPPaiPufZvXsD5smQJOfZ/JHO3I6sp7hicPO/0HB8ZnV4dgZq30z/6u
5BIVh4Q92R90Ve1xpZ8PWuaDUl2D6K9RLj5l8OQ+YdbP4xHLyfZqBRnLTyNDyezOqmGPzz5eNp4H
C7tZQn90LRAK5TMb9Wt4ITJycVqWgG9kMVjzc9vUa18EoNZ57Ebs7wwqHMel8Z8Jj8grkHwKwIfc
kKTLOicfJlWeSwpW+h/26QDrd6iKweKfSiqaxw4f3gjQTTe57YSMZNUQO6EJk8e52GRxYq9NXoHo
XntwVM11M9dafszPH4t5XJ3hxAuuApMEKZH6bYCtbXbO/uooQFtKWmR9R4qnCZdzfSb3MGyMOT7C
3MvcPkT8ScSaZVNju6XzqTt1HCBesAyNyxNBqBY67dSa1jb+aXb7/hE641+VFqCnk7iCwrgrYytw
LDgdXT+2NEsnNMhy1qinuaLUbg/6ecm/bW0RKifP7PLNTb0KKD5Ei4Wh/oJCm8gzhU2i7u3EFpti
t5+SexqHnZwuDnU09BrxcWaTio1owjEsBCz/eK00btx1IcqfjLA+3HSyCu8ROz4LHJnrItiWr8eE
KRU/RbkAaI1NmzS804bOqdZNJuUvRSTY2RQ6h+oFW0RGFW2UpbLmZPl0sTZO7MotGmpFxXqXiNxR
oAR4FQBjxUov3AumnNnPzHVWx63VLhEI9mFjL9oMFXlhYyl7aSS3HXXzU0Mbu3W8jXmqcrmNtnD5
J7OLlQQVnb2xJHd9pGLzsqLAK/FCZ/Vz6Hb299+pK5t+btHwd1F/fAw5hxBwdRHcjGVy4b0QI4x5
0fvchP5Chv9RJm58UdX8/KaqBTnDdSlUymUDCs92jkvBxUdArWlAcWB9VcT2ZeI5ZDNg4fz5f2S/
eF+pg8Of9yJ+8n0LCB9gjMbEsM9p6pZiF4S21GueaAWzlxQmPcCDTPqsRQ9YYcR50y0W9uJi8DOb
N9KXOtc5zzcnHsvQtXwK4eYEw8Yuc65ZParCRuD0pkOadQZwUrhLgtnooqi11GOaIlbe53Ara3Lq
mOxkKJWexBmNKRD9g4g9uDwF9fQAIzYnnhVENJT/hCH3TvhiVF9XbdzM0GYQF9stXCcDE2SnRV1C
oMgJLKawDxK+eoe99ylWZD5+aua5USKqjPBeR9W1MhZXYzPuO7J/GqYigN29PKOrFI3Fqygx2Jzu
bYrG5CC5nRq9Wi1GbFDoyLMTlo9r327KaouEH9xsLuQFaRKPRtdz542aHHHXSusigt6kxKbj6B95
blNwy209AJyH60rdJ9NU/nNRijM7NLkzzRBNcGOojl3q7G2jriZJeDGnyYKDp40t1d4aQTh88Bz5
os9qZD0TBQQMNZiFT6oI2gXEI4Yi2z3IoANoPnKpRiAlAyPAHBqRM6BTD0B7accKbBWW+KWHwp8w
XLREfsh6N8SLnJ1hGncRs60FLF8LhFkwsyhd5iJBTZS1YRl4jnVWZ60MYjNAYd+nL5nudc2ow7Pj
vQ91I+cBJIADEIGP5aWwvk6iRu1ZLyYCpbN1qM6XUaJUZHqJX1buJOVXBzfq3LJA4Zs96GqxAzP2
gUAXvbGwYgxXvSbEmjdqt75CWsgGL3KpvkI1K8GMy5RdhxKYbyNd8v6SiNp+lBrZ3RSJy6666YOw
KzjaajZgaHmZrg9GoggSXFk14GVLETLY1H4QMRVf56TX190tYVmrZWx+XUPkN/FPeeIliWhHlA09
N3FdpDlT1wMp2TdIIgM7Rj8xhrrX9WPt2ogNnN+I4Jxu7nxoV49XAS6lfZjTfmYZRPhlQuX2JAIA
zdpvyAYPT9/25VPGYAfTpjrYNDLVBqBWlqzwE2KXAYoCxCDQPCCw84NxlvMiINcOyJ+Y0G5nhS4f
uNBNjGFmZt6OEqEv3jqyky1o9VEZIdDiTWw/BOgxNlNwMVT5MA6/j2tzcGfhPb9Gsshvo1v8CGPk
6xOvGi1cxaVEviWE0O1J82BFxBOd2D2IxfrlPTN1VSM/noHbZaVCNtgPJ4iOKvmeSq0pSSYKYLAB
6atEFZJbTdkBIxHUFEZ7ljQYnRFrYQ6BiKJgOGBh59lbIhuBQ5E7kdC3ZJm4sQemX8k8rXHjkiLR
nVcN4CzW0LCis/16PE103UjQ4HuVlKKPLwhR32T2zm9SgmA2HAGRp9y2AWFMHmhUHnYm3LY3pCTe
1sRDZ0XVqV+X4AtD+luRy3tgdwGaHb87N0oe834Ze0piksk7wwSnFlQa6w2cz2f1/aTLiDAAGEKg
XjCmtEAS2u106DoR1IdJi6dM/L3ZSm3S0XXJEyHhrhKo0z3af2K2X/yzuWPAIIgbamEK+4NpJeU5
aPXZcBw+OjRmTJtj0Xnk1yzb4NAI3CxgwKeMYeO6uM7rS30VX2BLYnPiO6+zRoxglr3gu4BGn+Ji
iosEDnB4DxHgFeIDyGpo4u2pNdGuyH0L84kDAETtiQMwPf/gm5B+DdWsuUlZs6uyf4LN9+PSLXI+
1g5QqlGgDu+xA8vZsvqmFFNS0lygxz+Rm176muvu13zS8hs0ZyhMh+5lWKAnksVtj9zlvAEszjsl
Hti7AaUIY3LtX4lGS+pY0VUDLDytJI48mDikQVaTuJvcijLg451uoFXqAeNjXNBE8WG6+0+pdjsr
OfAW4lDEWM3XSP8HErbOeVa+ayIhaD+BVc43dpaROlOHbCXsjNO0/VwN4DhvPmzqdqADw5dVHSL3
3PVMeQbke0cD2sjGg7Ejb9JWLmdfoZI1FX3xNQj59AeOFuEgCraUVXZhF7+XCXlwHl09DdczP8ZI
lx/y+aypmi4+ni1ZrfiJF5WzwvJ14QcS/NYokDZA11UMjUlguYdb0/2llilSA1/QDHVf/PDtUdq+
P6iB05qsDlWNmkHLGNElpqw1EEGGUG+z8AVGNZLNqzwhkfv4kiXmDjNu7HMdZWpzh20po+uw78A2
bzSYqQkFozQFVvhGt3+JKxS0UYCIkeGm0OrM+veIQjPfIwobvVvxkW8ptFwQovhfuhQ+eouXfa8Y
tunoE3KmujF7zMZRx1G7V/ZqdzcWzjoSIWp/e+FlsXC58tI7Fxsz79oKnHj7szp1L7meof7Ucf/m
aN070NBEnC2tBnfT65y370tFCUadd6kENx9uhGxH7peFfu5ZmNabr/1GS8tYoAJZ5AlbYOVSeZpV
G1+trfD7lIDTO+WyaNJ3FVRm+psyejWtc8W2jkhn22+SrjxPtyyWAFzrb3VvKtl9Yc1rZmdfuCAk
DA24lEyQNx/OSN5JW6o1NEzBasBLmpB0DVlgFmGQARcGBT+G3BhtksGGWT7s09Z5IhZFsONuwH6h
huHa5amR873gMeeY8UiidtIq0c5CmJjCLs3SW0fjm0ZhqeNt+FfIqzN7i4OwunQJy5NDH6GbBimY
6F+ECU4CBk0SAfATHVM3C6AvgFxnPG2XzzkqXEB14FDT/iB1YvG3gAyh++T6ZeA9O8EGT5KFhvU6
STMLbBi2j2qsu5tK0zq/zIH2LaRaaGNiqp66A4lt+HWtJpKMtdTYZfFZR8qdnZ6X2BI06LrhULx9
KpvD1ynKx6w2wJ6ZkjYLy6RkSoWa3d9mnwMRDDdywTAPj0wpsqkqufg0w5MP6ArjnRVnN6lWI87r
mXFkE+KVhghboYT7r9EnZzJFTMGJ/hbEXeBfmSKONxFq1HVYTDvo4GQZfO5y9TRFYJkyEyeNmufG
vVU1C3XP5mimTskV7S0h4/dlYSL0yvr7am8CY96StnTCjmURgk3aWajJ6la3WOZXySG1y3HNq0kz
cGwNIAvoI182jfKixXw7/nJD4JqJqOM5sDa9lIPn22nT/7eHEpKLxFC9fiVBp6Pdmw8fb2rLJYFR
++wfGd4af/ZGfahBg4krVa0F+OalilkbpmlwtgXPIn50wTJu1RsSLQIojwXNkhanvGja2kr63YlM
A/PzL79JVJr6nIPEQtKLeAvSFF64xHlIQRFj8MBMzzF/SbzCYtZSCw465VC3K5jYx1gCvFHZx6YU
Xdj8ERuap2bhlGuSLLBxqE30APR8RsTKqGDz9KH4PtfyATfCDNYAhRatUkVgjrNLK+ZEk8AazdKU
HCVQn3fxM6uaDL4vMQuFwQLEiI7s02qbQJpue69iab2JPk+5vIZmlU6l6osFqfwxfL61O4STFOFv
iLFovrTNR6PaI1nmmU+JIkACA5EeAN9V/byODafWOVVsSKt9qSAjfoBYTBJwK2OYe1dJx8s4mbwn
qAs6HhA+kS6uKIEinUuK3ILFQGool76cGT46n1AZfeg2mKRn86GcyYqqbd/1nct+5IM54GZqPflX
QpuRWgO4XYGCkQD4vNk0zDF4MqZF/DfZnIWkKoOb0uqcpDWOM/3MQruzRgaTcChGk81zzi4qR+mi
5srgy0rOCDW/Qvjm2nw2xGG89YNDY2vquVNes1Zp/Ke/+2J//ss2/T+4Vjg+QrNW04ZI9TkjubiD
Ryng/hEhE56Jk+rFDbvndHRxCILGpqk0EzrVkofMM0LkowqvNSmoaNNoDJtzWzuG5fUaiiF/fF4v
t79Zdh26cruvlMLE4BpEbUx5jFLaWY4Yfnf4eXo0RIZ4KKReJ1O8AB+nQppSh06b9WxUeIojqsio
f9wd2oTYcEnJf/hpkcVpOExtkdbrg/zHeoDRalGQlZ8nbdL9cpcHbX+29aL4R9HJDTN4QJaKeo+r
nlOtVoP4dlScSj7QJKAZSgF56DIZFoUHMhTXR179+7IQtudlemjoaY6z5qX6MjYcCBjSO5wflnrr
1q7N9FMiFa1qBMThJPvVekEvJBNOSFu6u4F4OfKN1PkAE0CKrX9OPkU7v6qam2GJwUPMT1SCfL6d
aRifER8i0tn0qls3piiVSG7kHhGaSkkuAFOmP7wfg5Ho2h4Ty3q9m5pGtPtptpqw9uoxPfG5zyyF
WqdioPrM42QnEkufCqx5L712weXqwTsH0HpZpN5ALPGTaSgm+/4SKPbX1+QLNvza7eExV/jres1+
fu7YD4YRSLATUc3fWjWwpNuA4J92AXUsj1NkdzN9Hj1OfWsLic9QqJlGJVrYE0CvJr2jfxge9hMc
4LvF2s+VKLz21mFfDumEUGVtzw3xR/sX2SVXdOMVpNY9OIBKz9i7udpZtXQW8DQwAhW2ufBPVKFn
jbkoDgzyhdjqPqUhIsgeOwjmon0kNIRbbwUvU01wyrC/16/xyHezfH1tOAHL99VcJXi6XAUzBPMz
Lg7BbI8/h3/lD+DvYsOPo87BMOjlhH0vZ2PjKW/7qismY1+y7fE+rn5eMeYTybYZc/nKfQqamkwq
SQHPo5hKCbuT4K0fPYECtJ+s3EuoyQUu5zZfF0NOcOW44XoN6dzmtmzs0SiruER8yFEVpMwQK3Eh
gq+Nh3W5jOpLLf5xhOoRQtpMKilGkaB/H+VTrZAKl5NzFvfoBDSln2VhGP144eTPQHsL9WHJkUC2
fr5lmHaTK6Vxj/lUXM2MnJk5KQmbJcGUfo0dDRsfcBCNwQCNU//yJTK8YwtwMRd4FCAHwLybkDmZ
0IwFTnPpYKd+qmguZ85RbFR8Jj7JFY0/wKX082W3JkxScjyCr+hkfKnGswwYNIrkekcgPOQzklUX
jzq22cL1nx8b+0exPIIaafIYDXxz9d+CJDQpJel4CjWcJDPB7580OI3VEYb6AYBKENb4GunzFJGK
8paskr5b82xdIYpw7DEvh3RSrLQ5YQwNP/h+wlweGwpxrR/BpECDOB7Q5EYjwz/eDzFn6Jh2TBzk
Q/wKwIFD/Hvt7BPDAu8EdyVb8eRWSSkBIgT+rEA5JniVTKeMrcOkmD0OqRlSD+lQn4eiIfqUrKOa
/nxYqgyGFS1Ev1p1rvdenYFIjiw17kS2H1HFOflWzL164zz5rCNMCzHl9U0XiWihXqeUY9cBB3ta
COPiEgbrFHQBjyy3lkQ6oUuAMcoZa7avdrK0O2kwaDPe0spdEE/gd6EmReVIDtfofieQ7uYYgG+T
1E8N4ODlNAW8PMGjExCwGvG1HUkUd4wUlLLFXoRq8KbKnVig1wkkjFag5d8osPUOPTgOL6cIgesn
7TQBLzHb1xec0EZs/eNWrZTXPRTuf0huCEXL/+mK4eUMCVcHNQa7ArGKlCYzM4ovvp3b3PkiQj47
/X/xazgU9Gi42Z1wt5OGT9dhOaRsncdfcpwsVgTlt0SnyeUEU7VGVdUpia3aKNhWDaxNHNovWLlu
p8eqVjL0GZLRWFcaUD6p+UOL68OJb7QUPjaaZ0J1cG/oivZZgvXygeBsnkPpUP+zZCoomF9xpv0N
MMtPlaUMVZKy3vZ9aGbIIuHVDMOzxSLSSPoo+EwSZ03me8St23uPBVhQEvxCjWj+WmBMISV9oa0D
ME/nfUWqq/hjaLdQ68sNUKBNp6gcJVVKu4EHjw9TlKdG/Ce/TjJco1R7b0T/MC/tdpvHOecONCTc
uep1NOibTIRdFRHXF6upnggccZ09rcF96f6F9caLlhkuy9/Ze+rDCMLiywGaKNYh5IA+Efo8CKzz
fRPLdlSrPeiTzG69/aOpMZjsVaWeSP9uLm0cxEoOps9E//aTjocS4fy8uANuEZ6NYcBfvh8u+1tV
fZJa+Njq2HiaKZIp4Qgkl+RwChJ6JQRlXDCfSrJv4GSF9q78Ajlb6Pil23h0C4B8tzS1F/nQX2if
mRYGgsKc/EACpKRdRxGhv5QeIC6hxHHrn9Okw3M30bdMZCXhtRttnYZjfF0xSsXFTeDsgqSmCz5m
7TLyKyVLDt5yTh4MPXlPzyDr24oLORsI/HAM6oq7iSnqCdePzMiUUTjeqds8eQNWSb9NMRTbOUxO
iZHY4PZ8Np2a/AjpG/36CmK7+6E+aMdoe/icfnWaSmFxJmiYGgisvoM4Jwna5RwrmeDKtKuZladT
B+w4cy+IkyLeogjKAqlM9Mx896GHZTDMJoPn8lp2HfXMQzUmspXArXtf+hFLZsAq8tuIVb/daXg8
RBIKh2Ju3QDg+wupkx+ILbYYJMBHVvwljZ+ZGOtx9wE4qAI0FcKV7N1bSrR/jdYGuZthe9fwvUvc
jPTPYd2Hs72RopL/z++Lmsr7ZeCeuQy0GxepA0C/04D3+d1Y119eLywJ04plC9kqA0+/XdOhgUrP
8DmDbCBuaOfBXI04JrcAgSQHiyOb+1JigT9urK55BeyJRxblulypLayE6lUutlAhyHqPVJa0F9NU
Bum1Owtziqgn8P5jmKuDxEmxBxR2z0g+IWE24B/62O1B4T6n68sOZYPQ8wg7uwYDpZtANptRieUS
eGlbmULg9LrXHWLYzLwgrb7cCc/QBpJ3pWYmd3YYHe/sN6kaDIozDB3SzbpkH63Y3l6ps3MM8B2F
SnJhAg1P/gPhZj8cR9W7MHmaJLjslhDtsIEX33O3y+8U9JCkUev6cZm/aaEc1pKfdR4a9S2Rxa8v
n9RrDLuaJykoDpZK+yj2hy/+/jBf3YmjQdb+2/0T2VN6+tJBEL2cBaUVn1F8Th7RtE9TPAPNFu8X
6pRb7KIPdyVF5oB9JsX2hH1L2zcf1JQBgdTEFqk5oxrXY3scSpY2+8QtN31DE/3An1NtoHRxjf7g
pNAbHnKFbmMC+ATSB3pl0xV7KJsd5ceXVgTJHboWKpW6YGz6NH4+ZgrSuHIB3qrxVGMrBElFyMwU
B9NHK8kXfZHcVfoav40d3xQlHJfbQYrY39CrFYMAyaq7LHhGuklEcsw0jz2q7nvQEx2blAkNeomS
lj5HXHX8XMX5hjEKj5TCPN69+0DyumcsV+OQd1fBVFLoE1YRbtfWRsRYItbBVaX/s/mUaGqxGkhY
qW7PLuZpJCX+doIbLf3Pgr2fB/ws80KI+rwfatltcZZMG4vyuHRg+j1p75Tuo4x0R5EyUchVlINp
X5jpkuIL0twSg5tzpdfiTghEQx9kt009heKdBS+DVeECGFQcULbi62k200NWnb7yFrkAnAmXZ/2K
HYJi4tPILJv4TH4F9E3nyhfZhjhz2nJJDVl8rO5DbMmpSiIUCT+tIFCSucTTRUPbQqCDtKeZSPA0
lmPT2DUX9z0jECGqtlHij1FI0Eq4PLArLxT5tVWOwv779cKySusb3LZu2/zO/1kS2bR4LTyQlfgU
jOVwM9sy0ivdttnThfreOz8GT77s+vVtNRyd5xSV2gRumHuv2Fo6PuAov0jWSMDsJCJW1kSO47vh
R+Ap+0mSIqB794S5uJbQA3DRZhYtCCOJR5puP3lPOlkqByTeFVSno3q6yOzLitn2Veejm/DlWm5F
0E3e+yqFFobGzMSw1ZjmRqiF5fyCElJyuyfLYM3jAE1n/KUY8wyU4gsveWLybofYumRQgxWTrVAO
/gRJX9j/MprofElm6j7zsPMKLmYYUM8pXHiu2uXKQWyJm2HwDxO6U0Jmnn99Fzb8KS/NqKn5dMOl
gJ+xwuvdJWZCMGCV+POnRu4GlGWi/6nIHkGg9PSH6y5dlbKz6AM4uAaAMOsbRoB4gk6UShr/qQ5E
8LxDPsSq8ehinqkiVcGRhYvFY6hA2H2/tJYfJdSKvBN7uKRmOzNEgniCaXa1zL+R7h95viC+/kEo
Sg+6qL7qM41gLIz6hx16LyIRWzWjHa+1YV9Vxh4/R1q3gPSXMCczTQy86YTHFclXhURxcE8SGHmu
tNorhYs16MziLchwM1CHcdbV2JXzolL3Ys0W6GzLHH2hUUH1hBdGsQ+hyod9hGhzLNFX9FnGqpPq
gSCKKY/t+g0j7d5Umfk99CjKLCTvz4StY70186IDkt9vs5kS8Cp7yHl6+hbsnJWoGAoOUjn5GDut
Yafd4dTC+ZZ0EBlE7bVVycdhdUBILoJVGXxy9OgVlk0KbD0Ueo/fMYwRFhA3EqpzjqOzuueyIKb9
ldAx9DhRgcWw2EFx/PeP2Tf5Th3ziuhYW1yDSb0XHxbIB2fW4K9hh5dQFD8dyeVaci09YFvGglFz
abpflSx1dlQfkYwik4oqRvglVe/+t3uszQnqy/3idRPmZ+W5gYeUP+1ujYHAM7z5z3pL30fLM8aa
0/DOeq2sYL+gTOX/PsgFynBjjBMk80KyaRXlvOKZjkxSjZ9LUnTQXy8+pwoIn9fVaQG2NlGNy7TR
MmpqAnTisbdXACfg/ibZGB0iSx1ImDCse9S64U8VjR4joWdXDqrjhxfzyqANKN+SzVbn/VzX3vau
hbjQjaoceIBxeETy3yZpX764nqIhZpT3MQP4+Vb0+cBudDUaXc2OkvA9F/OO7Z/CWttQZ5Npy6AG
6pKA42THi0+xw8Qo19kbWASvs4PEjQBo7Bdw18EnhMHNL0wmrOc5VDRTciN5J60WYdCxCWdS87x8
AzcLxbaP8D9UYKyYGuvL3GtuDNLSYxj5/HzuANXPUxzXWA1j/mPu+dNrMCW1aXzj2bnMGZO010qZ
FSq8cXrMAeSDsPzSGumar8/+ZcZdCcgsz8VfIKaHruqSmAPnnqvfRJu34MPWfe/+4D6bJsKYds43
gKZs3Tz2o1hvJCrCBBdIkze6lTE8WxR5HOeas01XgBU+q4sCodU1lygdTLpoFYjQ5yMq5QtHlZ10
Qn4jnfiKXdF9Am09xf3C6o2nRPtOqUJjU0IIaPBywsujOvVAU/IVX6kxOVzpUM8xdkJVNnszqMor
0xYi9J91DIERNWr0MujFPdWe2/rUZpuUFf24AGoMwIscMAxz6UX5Q+g0kaRV7BsLT42w4L5CDJY3
39Zrpua2PCFXr7jbEyihKHiAVN3gM842Ipmkg6ZZfyAkYdRMZLiENUg7auiNmweL7ouaC98MBbZj
AGw/3WsXCISI8ItFxFnJYBF3t60U7ds/gf2+6XcgOkIFyEdoOEmBB3xmKPd/bZylRuUFz7ZZEZYF
mFsm0op/7iSGbOR2w8w8qF3wW26PV0kXGGqy2Jkto41+1UQ/l7E/ru1ehvhRpVvFbVJ123ZDI0/F
bpvV3NfHJWRGsOxmNP1SLOIvaY2nReG8cl6ago1Wab9Jq2IzuHN0ZT/U04Brue2iqEsFBQOFhLoh
lifYAHiGNYJ4wjWnAGnoa6eVrs1En3Z/31QC3bpvWCdEhtjVgxUCsSyaH+9zAhXMdWpiy0wI7HOM
sGOFAgaadWU8QAcExBjKcs3jGTV5qaAUcK5dFlJOUWjH5J6AN5z3pvLeTn2S9cb0Chq8W/Lw6NEP
ZyL9CWPnSnZWj7Fx+4XdeQphNH5oe6IHzs39/gX+CX/1z9gx2C9SO5q2WYxXsV9nUIIQP0FOdpl3
6uXb4oxuIo3pNrfjDIRAf9Bpd35Pl4eFWFD/gZt6T8hmgdx2T9HZl8MLSi9RwMPx8KJPut4jdavw
8Rz3jaLExPQAugcfClOZEQ0trlP2oum/m87EsOqTKo+yWbVDP25K9pzcW1lHclW14/EB+xnBY1Wo
vtATB6g64l1kIJqWMBdI8w6NmFgNxXWBQ7d4u5hNEEA/TAcfTw/EL27UzqXaMtiF26CKELcn/DHE
isRkjYLEoX69pon527mCgAD1VwEGC8plqWJknQBB2XxrzESG+NDf/e8EH8sDzrPcNv3z+G55tZDB
dbAcwZrnpgEqnaSGaQq3Hogsm1fjkZtfvrvygErt9T7JQFXL3ZO3tw3Me4cYqGTLLmoYo8Mo232O
UNqWTwe3UWncNVxr8YU3Y5ptTR7zEVMK71weyFnPud4WMx8FzC1N1V3VyHTRiRLNwsrM0X4x77Bo
sjN13HRTWwg0D3cRvUsNVafvb8fz7OD9xhDmrbfaIcCr0BnoAq57Qsm4s+gopFoI32J2lQzAERON
DsRefXHaThhRD4nFJdFeObUikwDBgOgMWFJNx4iSesZbQKto0Otvny09kVQgMNIeN3U0x4E7F7b/
ruCouaz9f1+zgoxtbbin9xR1IBg4chdHxTRR+FgEqi1urpIxuZ8Wxp9u4I2hTpUnpmr7nlJluxYO
8MvPdpw3u/E9xloMS7UHmm65jMZ2/Apts9a231QdBPTi8w2AiqmqMGdmaJBV0M7keo7EuVAUL1y3
TtL7jmYBpNn/ljL03EADaMNU0lH5lkx7pxJuWChbwl4ukqf3r2d4O1+rcV+J+WvczUOFMp5GxI2F
9ijpgukfnQVMnErJlIRplmERUGlLY5WvbjIo7DdNPeI03IeyAoKHHm/IeJXhP6kXL0cBQVAtEDBP
4uJuyEMT51By8xmkqsGlHJLCpa0d00VVQpFiNFOqxOv9Vn9X1kFcwaBUfCmiLxW/ordfy/7ab8KY
k/X8iUnKBaRULfIKcAOEUsWTxxgaPSP0EW1F2BTE5lVEinBHUKQ4SAj9H3sQxNLMgg5ua511JJTZ
NSxQ+u1GIlXfi+n2W5ggZkk55hN7m7WFFnhhl4sN6WqqKbAyD9xKtZOh7n822dVcmDf4X2B29li+
kFooTElYZsukfO2tO3F9/bqzfYH/8Uw4GS9FxR0xbIrS2YHZita0LLxUm5yRc3zfGVDnZFysPV1Z
G1iwDi1jIem/kxeUuRPYoRDB7D3xnpBvq/vjwClQQ3W+S9ge0C41Qm99cNuWjG6o+ducY6IASk3F
SnCM6mB9068OVDL9WNb6tudxEtqEvHimZiKilq4298UTadNAik5lM1C+wyH2sxAzveQyFnMd+930
zbKk5PQWb1+u33IwPdTEemeFu8+QTXMhlUdpeH3HaROC2xNS1eioqcAJgNFPZi01l7Aqq8XJ305V
0KymE/RE785ZSzXVCVfLZFSQcsuABlyJ1W9CuzqTBxbO4a05G9UU9qqPgBlzAXvUExtQ+BBQUHcD
ymOsXDvszIckDAWVwNkPSHkbyXhHYDSgz5wXskNIdl3uU6KMbQ3I6q0xEaIa/AmG+o5Ub/C6ooVS
XdaS8S7+AMHL9ISI/mJX29yqCju85PHyahN5m1cxcZRmMthwLF3lmFHft8Z692+YIx+elKzae2Tq
hDkfzXTHGv6/fJqz7uJ4Chi0enq44z37O5QksbMqdjs5dPP2q3Bs5Mma2IhK1fMoMGSh2+iO6AaF
BGoPJn4fq2tN17Zvd+2TxvdoRR9oJ5JRTmU5hxgJmISY/wyl2eCjwosabU/0jzUZ9JbVwrFJawSx
szvrg5bA5dWab0ZbcypvI/zjHSTc8JeFiTZsiEMNbl5zvifqOcPLIadxq+FM/HwYa4ziKXwRxX0Z
usyr3E1RlzrtAX/W5hZPC9AuhW3CzFSMrParXog8tRO/4mmrSiOYN+3ZggFyWpGVASdMrG3Dgji4
HFAMBselRvtmqNljM7JWXy26rX+hmk2HjjpPgRscdcK2czBdW8j6lZlJEH/6cBxaoYPCnkt3OTUV
zGYJRq+73kIWmnOzegC/9xvlmg4rTxrFti3I2sqlx9bs66ROoneUV4aYWDstPKRmnyvNmlcufbVB
s50sSbN+s3+6OcJ91e6RgnKoOWEjfSUZvzgIgu9p5wHJmsY+ub++Eo9uWPl/apl9giht8Zsjzr0v
hb76Am/vDT1YhwcrE5hcQh1/DuTT6HsnSgeFGCWKadZCBzYZC9ANqiAIkt1bx7A4HNjOdEC4LdbF
i2ywdQQr16glYlxnSQdJfZMk59cKr9FJinNUCWy6cged9X6kT2emz31OB92aHqXfCoVi17tBGdtk
xMw8qF3SWI4WQXZGJlBgnmAsJhzCHY1BlrdCnTau8/3og+HTMY8FaGI4g/ea/tKO8lvdz99dqLGy
ajKvua7B2Y5KnuqxMyRhXaxpgg26dTNEDylz/eLK/IWNY7pgIVXafNw4LtiD1WDterTpa3iu4Amz
icNHOwRZQcyBWB7qK+X1HSAjFXCP03UGthHfara8Xq+FBxqxi2WShl02yi3/Nug/yVkSNq8WcN+u
uCzlGorU9RwGAfYt29f7JzcE8NOOTOX1/DwEOh7gx8Sfz3DAivlUskux1rguyn/E/bOp1tAXodRB
cEkvjRKHrQOZTkHnfNpGZDKaOX9R30V1KJOGOjgrdjZd6I0DoPshl1TMhZzaHDLCYEO8pPZAOpMy
d7+en70gXhY6FAvW7XpGhqVHp/fayqlVcgsqDbVWmsG2Q/hWS/l4H90XFUETG9Kt6tiB2o8qPME6
37duPAU7YqTaorMVXye/nKs73wEY1YL1zy0FTvXArG3kl0m7R6ZBWl19WNlIDikn6yFNROhlNWbM
nJQppDqYwpMN9l3VIBf8XvemmC57sUguZXleJI0XNwemtNYlwsgAudhF3Zcmh4+JkQ2NozMWwPXf
uXfB5FskpO1HJ5k0PRw0HYGTsQCI8QkHCvK2WnHPv2wbvaBKZ5Ru2aQsxLql6hy9Tcat9l9t8inR
pz5DAS4riV5J6GSyP65cx73PFd7atPHSm2Od/Zio+j+8iXUTkg55NqDXjwnyDHTNb5I93rTvT22V
XmRAyoGR72hi1kLVO3gJOGpC+Im6b2azAlfM4ZUZctoirzgy8Y3Lce5YXBFLzVNVSM7GSH6Mhkfk
KF+jMqHhbPawfM4AaZ/3UBEIS+X/myGrqp+il/+3qvN8vnzakALX0kcxv/TYw134e+3ZrDukYPGL
Vv6q+/8nZCVPhMumKHQ+hFvmjVhG/+Ty/o25SxFSODzuT2VjvKqiVbJ4s4zOX7RnZV1bdqew3gah
bEI2zvWaMqJVWf55EjCBZx7LhMmqjBP+CCV5WtEojMbfTTcGv5GTdQ1UwI6dPRF0jbroWxGhbAN8
Nr0JnnPWxVj5SY441ETQQnX3wd/Dflgxj02TZCZIEsc7GWD5Z7+twU8oDNvlYNlN05VnIY6I+LxL
J0B645/f9BrREus1zW9PXRc6360LJvs/bRUwhbJ+p39LWouUeCqMwmyf5ZamyjCzJrUHTL6txBD7
XAyqDmZUg4T2hnUFHUD1Y78WqCQedFJGC08kqYrbZ7gxbFIQN3/IxmhGybzyu6CCkK4KzLBw7wpA
92WXw9TB++RNCfUXaBvKjZvhfkEBtcxtjJMmtaVhG0zWIMcaTgdqXAHJNioRyKtQN69PfPAsa+qF
kvjYi6C3fsXwlEXkodV1jrstLegxaLvoO0Sv2GpeGN6Rvn0jgxy2UopTbgSKlpqWWERDXP/Z0h3+
qWyl4fK0AsnkpkBJE8MCSM2w7W0LLqU31pcKKGd/5Tp27hxWMr06enXEsYRVI+WRWRjbdIC1B1NI
TE1iATTUCD+OiZAtyEF0S6hRJQ5x8K54hjDBMCK5XYv1ggsYcWiIpkGLjvcRnrGwyXCQU6elKXQQ
2tggo9Py5ZbfWZk7jWCU90q6271uf1hmY4vN/SraoNYxO80W5nF/3d0959H7TJWBRXvZilWK7oFw
YicAjQNFVVhw7BAn3r1noPK+YS4x+ll2ppZQN1Gq1k2wErNi5QE8M2JXIhJ9ebc2ThYhGg3ndREP
R30bvYOtJA0kzIoZ1koS5CSFog60ikiD3fQJw96HK6hLUnWE8OB+leSbvoCupxHP7bnQRd9ibjSN
ZnvAiuJEbV10jY4DhDCaj6c5K6rs5LTXsJIp/AHhR5LDl9QVUKYIPvQ2XrsJaXsrGyoMYKUy77u/
OKxAM8piPRxyNLAUuNOS6k59kxO6FfJN/MZuQgsYEmPYgJEwIGRM2z4JZzRUR6BKKXGi+rrMj9iR
3rfjTE0nKLGNvrQqvD9gYTvz2d8OIlLHO9jjFZT7ZPtvlAOAHZXJ6ll6eloHSZgQbLP9WStwiS92
tK7UmFBvQ3pdMIFlciRTSTYOlXh8xNQqNJBunubpf2r4h/skv5eghkdf6/4GOgz8PqcUn0AOrYBD
LnZuQ0gNVuKx2cN0ymmPP6vVo3W94ytpIWmz1/KBRLuqocYsfI57mg0aeYWD59Dn1ttdatu2rbxB
S9dyE0dxIRcC1Rbtoc3Ut6YwHDpHiMYuNmA+gNPKFoGGoFBGZ2hhi6P1mwqkQt1/7rzrGxniyRTH
5+yYU7W+tAmq0oUjPCzGN+o/SIJZXIRlzdn4rgNBvZ31A/QJI7SIZtTrtnVh99Fj/E3QaCMz1m7C
u/IGdPWqrrFk7kobH5DbbS+cryx40gcf6zIzaBjpvpGs3DwOD4zpKIVbdh5loUvyRZKnOnMBx18Z
FDCwbY6+L7ZauXWM3TN+44bFnzlSeKyDlmggLuHRmmoQqSJfd/DP39xj4Cr9UttiYs+HBz4Mv34u
PIKwHJzzXfBwgkJG3sku9H1nnbgJin3rogx47Qm/OKaUudhT1wcl8m8fDLoYPsCIFz0WagQzRPsa
CJ3fIeZkN7aOvlJ+I8GMjQZakUJC7pNDUW7MvTcf4quwrRW3iuY5fZrYPJhMw8XYe8OitPbnjJM+
hkFY3vlP56j6m7JLY92JPQmjBY8UjLYd5zctkqwX86fb/b1gOZpAzkerGZpdVrdqS4HGcxAE+Dtq
x4jdB4HV6/T+wnaOoiIPM5okEkQmj8VICeXx4XB0o17fVF/CesjTtiSGBXwOqpw2mbYb/oAVK9UD
aaGyLxOaskO+YVfRMcVvEFkcYkzEU3EDR4j9YlLtl7l34oVcOWg2UlXmISzd+QLnYiwAcZ1/O7mc
gQNqXV4xMAaria2pb7oCwzAQxb05wvnLYO/xMx+tZknr+1WGUhPFJwiGwvkOTU+Tj4m0T10bbUv6
lmt8PyCWNnOySS04qIyvOqhmY+LIZB7a6BkYqqk9rngZxyo6BMhpkE31oFmFwrLY0wdoM7D52FCK
OTnSIATiQS5Ux5XIHS7KHGKd1FXr4XwPoLbe9U8hTaw12x49rEdyjVZ8wnIjDfQZ82VDHCPB0M81
5yQ79PhZXYke61+ICn5n/fvIccmdkVNWNzvsbA+pbgcHznEFxjA9E3AZ12acuYOgazAGIWodNl5R
sMK2jUIJDodnrv5alxNABIC4UgFl4BMOyzhwMdY+OOYFre9PtOVTDN9tBlmusIhny54qcvOgwLmi
k0DdxXBrlDIUcjWMVCq9tbtt67KYJpBWdxf30TdNEvUXkuTzTZDiEfVmXtqLxeDM150ePH+0KtiD
ytUULG0BFqZb/wfQVwWmxEs34XbM6Dx1EAAoaMusAbYrbkod4lbuw/Md31HMAFuwvDOrAWYaqDz4
gAwq1XYS/TIBfCgNr5zTSj1rqUrjH+O+plHn2EvhtuAqyQFVHtVXs8a6dC6A656/ZPXHM2WQ4UV2
8PKeLYzvZ/0fCIKto4gga5Z6hEUhg+E38k4DpUvWBDwiHCfe9A7JmDSGFfXzHvudLsyXngzCgc31
Nk9blTvsD0BrlYRS4nuZo9DiupkFEl56QwbrbY7kZ3CRm9n66Ik5y9ioTRAdBM/8u6XZnqnXuIue
MsimwPgkeJ78MmrIguWf0bFK5MMLd0KWZO6Ou8HBbDKOVP5LgZMRFl41XjizjTRQkJ40AvsCxbeo
u/+civuCxqjZtjlSbpK+EFWBCIwdeDh86T1iXA3R1L86O3NKxMXVlldtK3lPiar+WYeHzfNITCFn
wSORnDJ1XcNgcimgHjerj0RJuDcHNlUF7ALwSCCesq0M7A5rWNtvoumoV0znXaVPutEyGR3iJp1N
lSb5CN8oY224/w3moVIAsNAsjwyaVAwJD4HWEcXYXEkGJ/D0bej4IljguaIWf828VXkuULEgztNI
amrsoG7NVqyEhPn6KlFMr7MReQpM63x4jWliYtr6Sg2zxppbju7b+Y+6SYpKl0B4JW1aAi/6mREi
mPUfLQSd9VidfRjBbaoUoza3GCJuMGWDYAcfCcUqS0eYS/oH7VBtxozEE51Q0v5Nb0geaCz58RCy
a5+1YTCXLZiKO5Rw0nMipB/lxsrB62+lYkcpt+nlMO4qQ/H8tLTZ3kKcQxmIoqne0sLUeURVE1bX
5X0kSlVYbR+4JINbPi8ULI6g5y1xz3s81YAqNviFSH0usITO7lBIY1iEvB4VSI9kIb609XMDeBXe
u7177NPaY4dSgSAbQQ5m15JJcqTT9U9RLfBZWPMqXkw9BoJJhro+HKuCSwTgsq5lC+WNPz9u7HD7
V4IgZyzgee7V/TSc3j9qFcPa0Ad5e5czE4nXG9M22nZIeECPpAO6TXAH2z+z5FlwBZWqH5BuCYcZ
mSM7Dvz7qULTz7TfTOauEBDwqAoiE92QJ0nfqfyO8VwfLvmZKeECHj6WfayfAH1IZweNq/eXvcB3
mzh2jvVYubA3TO8btUQBws/+Uj6gNoPrflni2sZ/8j13AdIquPD0aCh1hQtyy9nq6lViZ9AcZ6tq
09RvyUvAqVfbSjK482Se2VhyZBWEu6Bw/2xGnTqp/3gokCtoUeHOep7soL0bEdvC5X+yleLemlIq
ayUAOiiTj2NbBKABVLRPvLp79MGuALo7xTQgNlniMTey+xWleoafM3nXImgm26ZJOLPKPmgiNqMu
9U9Ke8d9QT0AXFiYdMyp8co4nbVnjFyGLw7lfy3/4culeFn962Zk4lE/v2OvOlK6PHEsEY99Hhha
eMpbHi1WI6VnioeymchPRpgizmR7zN7RHxpWYmKR6JfuvkxWsNtxBWl1h4/YAs55yVYRXmZQ7m+H
vzuAADV4/aPz7mSsEWxsqoYaR/R45BSfcJj50thOeOMUu625njDWd3HVnNfrQhonedOa0ILiK2MG
cyB0ZMGOjgGJ4R1bfsHJePw8jI7khAp1W849iWc48OPbcCOSHfrO1i8lw50+RmfDBH+PJwuGsKUi
wlmeUR9d6WfnnfcAp1WuHT+/sxaVfYom5NLdc7vd+EfdzfgLClTcvUPFQEKl8Mard3UHg4nHxb6u
gaG542qN3eK1eT5AI8gbJdvWsDwpsJZ/ibJzXJmuTO5VMS9+F9gQnhcU6kfipu+mTewGEXO7/zGf
DHGIjb6YvZw6/L/TIZPupOga00bxtY9X7uhcvUSJi7Qnnw4o1Tt8/WnuXXKRRWDM24o1sSET23EZ
FJIB6cj4IlwVJ8i0P0QUnfLB7yH/Yen0Rw+UUH32UXSn0BgmW+LJ9NNiLjLv05bhtNkVJ9v8fKQr
3AQJ00pmEURWDmJO6pQctqyBlreEitw4XyzxAKqfp1/XTieqRMJ7af7G6CxvfY/r4RwvRl51dS6k
eklUnCzLQpTAHq009MUu5/ELehwhKOD39KGrfdkSzTdPDAJenRgp8ZQJHe3kqZdUdc8AjgQqyI5i
yHolU+TRs2Dwq0AwUfSQPu6BVQhQEeBl/xvRR1CPQxPopF/QkCzOF95CgB/fumtvpCf7vS7bHU5M
qcdJsQz8pACzAY+WcVkNiGHDbE1iRKKHjmaIxwvq9GK34XpA6DHSGwt8pHC+Sh3f4C5KWlBV+k82
Pktd1QZQ1qmbq7daIwddXBGg7ZJM+bzCtEIlLFHg7xAQ0mslVItXyNdNYQtcKk1RJEhE9rJ6uBpG
hUN0BuRp6Q8aF43FP7RxIbh7IxVLAKMRkKX11yeGoVFdweHy9UnQ713lZJ6PG7u0QjA2rtkj4X2Z
FzSqDZIj4mFxS3bADE8UuFdVYM8WBSvjXWZwjA5FpHpK352gXO+pPvrGWddEhk6oZPZyeCgpy8Ew
MBHJ9YfAb0QtlFYOIXab0t021XoshKDo1P3UFntGYBekWxudRYavVtLpXc4VNRJDbjEtBpSMkQeX
p4SlNFULTpN621J/OSlteJqNVEP5pMKktAofvVr7Sp59kK7FJtxj5khwo/sYKmSYSMLfyUIBCxss
21xkRLbUINmhmB/fmwuwcwaky3GtELEnekDZ06QcMOKsNAQggE6uCnVudEPtmaiUxNlW+AIaWMu2
zjf7xQPAyvP3bzhLM5B6adDcLbqNWPJxQPgQs9mESq7TILIHXBDsXRUoGz1Bu3csTnU6ONfS9m8C
FJsBR4wyCZERjJa1Fo9jWYp2u2pXA5rA8B1vuTOj8I92TW7pDMHFMYkIgiyccV8Tsw0z6sh9Vkrm
u1KoAMETxTqSu6SRNVjANPDOt7UBfrR3GzwfKfnIBEJPjF78y1TiDP+FoWXvFcwVg0a9BtHtbNbJ
wi4fI06pHooYDtlMX0EeV4ZW5b7AL6dzF/D3+KBVhecHfU5NdgT79pYm1t59szcpN7+crvw0AL0K
85d0QVriEPmLb90wOGVq6P10aKMAK1UXHzVqnkKUKkPodryC0sfQT9yEa96Sg98xbel1GhnLak9r
G199GLbDegmqon3ymtN/sCVILXDMl1JGH3inJfDxnWlHDxa6fH6NYMEJFk8vbwob+DXYeXNMilzL
lEeU68116aSc1DmqdbwmbWAJb66lH0y9VSvoL4ROqHnCVA7zGBW03bVRJDLZphq5lsfvCFwvCzU3
fyUXbLa54LPh9c1r6CY/yBfgIqXTPvV73hDm1ci2AYJdREh3Jqx2dZefNkJizDF53CzpMMESdN/L
jMpHicphN5hBwVHJNub9Ghm0q6Ov7l7wvY14ExwplEyw/FzWGSq0EyCqcX+CXL/NiuHtCb59jnm7
ozMyPQqFCf/WvlUYz6qIuzAB/cY0EFFfiMN9R3dYMwoZwzGAtjnSB+NiUDpWkYSqld3Fdwn3z+Ym
zEvR0ZjPrTc7nR7PtYBIigM9t32bgsw0tbFR2TX6QvFIOh4G0HHeIdb48PzhyoDYaksrtxdjHZ91
z3OcbOERc6dAw8gsbfbu3NOsJlrNF3IJTKxjbXUqeb9MdkSaZhqC6IC1tTESg0Qe/avwbWeGCIhB
6fS0k9BSQasiz7BFa65XgDlYL5jEF8egsY+y+5+3BZ1/q1x1uiDGViK3M+5kVp1W/j14yj2+ujq0
3AUiIbFhaw8/ApjHHtztySSOqSvMMVTkfPsVb13zl8vMXvcehXrT41WHow80+yI42PjwoYH8LNc4
aNg2WgmSYlAIF5O1QUa8Qs5jy2mKhxQ1c+K6tyHWMDd3K9fKEe9bc+WFQx1a7W66BaCK+i6EqIkl
SJ3ZSR6Xun5CG29qCzCeqHZ/pv0VtX6ao4XwyEUOoQInOR+JWhK9Rut+/2T6h2OcXD3fkP2jEtjw
6DA3xngBcIwum2ZDfKCQegZRVT7nzYwDEmM8QZNXx5MpDMYkTUek975uyM7yCdXWGTzZxmiieRkS
ZcjLRXeOEtTtVPuga/LTghrpalYniucZlDNKb0QzYU1/64MRRZslEAYXJkurOL1LIGPQNmlv40Mj
BKp0zV0wX6DQwxxRbC9qMwLB+bpiPElUp/u7TyxmMo2w9SHXCkwpgV1HOqiTCIYHcqE86uF6iM/b
+RbYBA/MKaUYz282TzJP6c5t4D9uqoKv6HeATE8ROybKoWBOF1XAiYKjJFqbq71Nr7P9xvZbk3bJ
YeEE9uCnufOAkm1XoRNcWEB+9ckd1tjA/U04udELvzCn1ht4B4pptEBAhHvIDLSjG/U5dF6681hz
5Tey5ikWbLE48qgDo9G+1/vo5pl4wqCidnEcu5oS+Nt0czADHgV48ixYA5FVNPuEUQKrAgQ0KG3H
F1yNdck40PeL+2i7Dtoq7fnZj94tTQizzMoAQuFMftbuG96rja/PfS+t8LIWiOJ0M81FvMq9u+Fy
qwmQlWjptIw6DYekt4hbm0dYJtuDggswVCWk7HA2HsLkEWSC+XTLqKZiIncbeY9PAVXiqu4+mfey
UnkFXBcS43IRWsf/FnBV3Q++d0ItJgE+v7Avew0JZE8QdjGtwN9rN9vDuZSAsMjtIsfGfDj3xV/5
+2Jn44+J7EgRu81ug6WpBGkeaAWmLWB2wtZ13eynv5us29twzfuSCn2ljkd5GFLJ+AXvt9D1hoMl
zuZ6rKoZHeLgfbUHaM8OOydEzS+szFmxe3mm+u7tpaywglav3OQZebBvYAZ1pNdDgDVxy418ZULO
RlLASHsdyhlHNrmtIUwsqWkip/9cBrIUYzmYAfEEyglt7Bh9HAyuzqQwjfw5Fp6LYG3dJrzfP7HF
sDw9OU5gRTeBBDu/IdoM5w7yXjU1o+gqUnoUDssz+m9Xfo9YBG19nysJq4YKplzXBxk4POlbrZol
KhDxmMp2n32HiOhLeB69mcLqtZM42ipuvHmjeezgTOluRpQcfz2Cpx+2p630nItlFlQu2AHwbgTN
9vkqgS4mOU8/uRdzpW6z/tse7NAngWsyCG558NWsnAIP+24mPYYPqEZpcTYt1KilklbkwZ9rgMpb
wZmIBJRIDRDFCs1BiGBKWjkILTNy+HHxBQq1MS2VYy00bLH1iOuiPjizJ3lzDX4VZWgiAD010s8U
0AuB+eJaASL5IPxYlE+KSdFT4iTQt/pFRDYXSv0qaZsbDjeEz4AgyWQTKWgkFvFSOhiQwPg9mglF
WxbD+w2QsRiMcGkmKMm50Vp9y2dyp26Eai3eJAGh8dEgN6qAiM4cF7EPCseqvIjjIuORRDxsDuiL
SD50BtPsitYCf7IzT2HCh1z6cZ1lqYCaCGsYALUYpI3ee83OpX/qnlf4TqiqJyDDUZ5OIjvxrOjR
pngm3WyXNl1GyxkSn5gjHMUlygw2rLpbwCPfM7jABDFryfevOo0N0Wk8h2D3l/7jJpsouCx7wXfh
2tuvk7dXg9q+OY1WmnXxXCSJ8A4Ps2GNIDR+5SFabzNkNmN3HT+T5/Elhfp0jb+i7Tp+s4lRnsjP
hxRQ+6PPmnVWHmKL3fbdp4BRGo4pY1dcFnpVrRSaUTVobrLUuaw/Rw9A4crEUN7+3TyoIc6aOgNy
ZvU7JivAvluwLBSI7NrtYhLu7prIlv6QkYCvg8nYdmFH52ZoBxWM8hM1BTDSU3nvMGfhKFNEZeF+
4Pyv/RlL0CCKTsG2D+KfwdMkf4nThdK11JRNdBtoZG+aHa2rik5lvt9FmGNZ/ye9v/8nrOnthukr
MbYMuqyy5Tk4ektP10OIGl5CnY+2boqC/RFaN0wxeJxJWlN9BJzoarjtzZpjQgKcvqqBURM1uI5U
UADW1qV/M/TVbA3DOIMHmI1SEiKPw6B+s2EKxfsEHeOMv7g8VtLEfc4ntR9vxChNvJvs2eRrjJy2
GJSPj+Lmy58iH9YXsInsputgZ0/Lh3zdgGeWmys2rfv+hHFCIyWKHKfMEapsaP3zsLSpOSCJwepC
8jwgnOHrVTe0t4bTFIC91qOzsMIauSMp+dN60TZDzhKqXblVQy1m4/hYmVg6JMRRmB+9I39SJUIC
ZMxSK1U+hTMW6g7ZFeWvQGUZAgZeaNtJa0iSdfZJe9uGB05ebs4PYQcBk/bgdFnR2EV3BaLyNhWI
1MgXnsvmLwgtnXX2XJiGW/yfXP1vOkuU9iV9E6pooL2Qfy7eNDd9HL+GUuMe/Af3s17HhSuJlKIf
3qKPiEqFSAGPV3ZNMG2+pnhHR6wJJN/nwJlaOf0JjKkTbp3eIM7ZoQLOfWs16O52F4zxF8wkQ3RI
CwvknLKjb2utEXwvx77Yc5Xy9ttqVibtpPBFVk2t8NMdPb18mdl8NQPaJyHmdPp2O2qu5cnLZjSS
g+PWGwBj8YrN5zxNl0VdIzN764p+w2orRyA04dF/+1YsGlvAbJTCONEx1stHcIOvxvNRoKy4jvg0
OLgohhfT02NMjMqQG74661DPbPpk7jOnBKIzh15QUD9bEwodrwQUVi04AVARx/OYjCv/d9sTe4Oc
N70w52rfkYqJ8R3zy5LYNS8smmUoXIdmzC7OzNYbsjeCSgkLvRmDmsWzIuTWwBB9tifzTgY99R08
5YtHznP38JcfEVMF9Ka7vw/kuIUNVpIf7esrZZ1Y3ef473VvnUHZK7HX0+O+qTeUEy+jR7hp3kwf
GTTB9q+G2f23+7iniK0WvKvovTS+5gJ6OODriY+5jfP4EfKrMIF2oDrvFyturvcUGk2qq+MZDwLb
iovded66HD4xS/C+Q9TzXpz3RbtzEWr5QX2Cmy518zjdBqimfvAB/708CCdjuacbqC4Qfn2FXLbm
xrESBgnkMKy9AMV7dDNueyVrtVgZ9NA1QofbpcKNbVh4Ze22fq+deLRvpxnYyOofpMTwWsQLCn8J
Inhf9qeDIw4LHgKPs/q5ZXfednAd7qdmuBpAdDKIKECUPdynYXk1w/AVUmukgkGEItDnBNYMiD6c
JYfFyObwHJt2tpHDPRZgyBleoJJTA4JqWCJA1NIq3JGadvE0y7S761jHKoU7abt8NzwlWIBl4jKy
i6xvZUeqHJnQoGzNWsq8PycoAb+Fhc5+sLyBaeDbU8s6OfOd/5WrluHz8Q87x90mYqoFhoAVzT5Q
Zmpa3lqH6ejVfueHrlMLBlSL2xH+iy946M682jH6L491rtHvGXJW0wSMCVj0FRph7rW4zwn8fdZ/
H7tDmqpS3QFB6RuWAlZPleNrD4fzDyY++Q+biPN8y29gamFpO9Sp9dKv5ILbwQXiAXYe5P9IUwn6
FVYv+eJ/xncS5tKlsG479Mg8+nbKTPkG+3lQPH2qkVUvd9XGbx881niXrE9A9DG9/IA8cMok9oW1
3A1i4VU08IGwq7x7rh+qAXpduOeoJakhcwKDaC7c7VP+moKlrre3tVVkGE3fTM+mWgl2qZ6/+tpp
RzvKzT41CVS4C7hCfE2XZWEE3Xp/tN6oH+RY5budlaMBuMQy+NFkCF/ysX1iyom8yRGK8JT6KIVZ
IFx1OnMKwAQthj8YvggDztaLEX47vb5xdRjLaAdxoH5ofMB21uS0iFRjcbQCrU/NYEH/lwvKXDQt
pHeDbHkIGqt/gyDmiWQPpTDIJzPAIOBwenyCcBCZnj7ZIwIBDLMWryzoMej6DlsprqtCbThhtrvr
zUDBqrcV8btpd4KrB+2Hj3yIPvVcgfQUc8one2fAPKXIjkW7vHYZr6g36FMOlY7n/CIRLhqDWFQG
Ax1Oj6ZbUhUYKF2vdZcZpaKgdvcyeoE2l3jfpJ8Xi975JtCyZzG0xQ+alQ6ZfiMMaXBAKiin99WX
gm8HbIg7C5vbT/pV0UUK7+FNM1cM3kSEZ0T6YiaES3rg2RPu5urdWI/OENVCu1O54YDMbESWDy4E
vmoccZI9/rFz6ogxp+m4T4t1CP+ib+YoQ4kRUSoMwS6zQ5P9IUnTcrS9qWWNuUtPVrcy1cUThuEE
nAbIRKnqCN/JNT2FBI06/GZaQ+SXxGNW+bahVtKe1x5k3yiRNWmV1CPC1oliUyR+cWFCa9o/rnHr
r2VDE+EuKVtMSkvT8wAvADEqdRh426Uhq9TT2oWr+Vbh91D19PoVmcdphJhyuCRzdnIrX2o1RMTx
vFINrvFSBN1DF72jugn8HwhlXuUqcMDtieOZHDnk/C7Do72Z74kHKa7BmFffvssdUZwIygjovX8T
FeAoKkwh5hpplfDXW75kbOCGOwvLID/OTiJUVai+ckO2QkC/LK5fz01y6xVXPp3I23Rl5dP743qw
ksBXI7FucEUj89gad4E+b6Zw8IwxGx6EvVKvw+VTBUm1Feb8HcRvBbbin536VCJqzTgnJSryX8e3
EEIjghMG+T/O+4X0VPjDAU1Qrv2E4Nr1ALo4yw/pxbnjtlSrBMhZk90o47dWmX5tW2Q/7102SUxW
Qs3ypn9LOzJl+JkwRa2wukTOH5dGVShw9+c67y/vI8bQrxcPHqHFLfE6SjQkFNG6SY9sfwBKhhyM
qBKsu3dsSdLwbHiLkfuXaeukV23xXOwXQPfua+frOCtFoc0mwZV2vMc1ly5/kaaVCF9uoMxDLlGI
lzIHjKredj30k4aF5QmnnmTMAUFQRwVaAkDXqxUAWsrfBTPh+YAdQqBcjziZhezER1INiLvSMfVs
1eRpgr9t9BfF/jJWDw87oTFtHChoWxux8MXtZV0kdjDFFYovSFJv373wL54io/bXuAQ9bcDHsla8
fxQVM/Ib2DcHlzSmp7p4/tgnRbbxUa1zMepvupGvJg2l2gQsGunUIaKwHVqiJVUm5o+R2+tRow6e
hn72UjqrAIhASlgXyzVf2gjb55g6psPk7U8s2JHEfgNkSpmfi0eUwIZ6ZIRxdZwMcQy3fXdoiJH9
Zi+8wlrRZAd7a2LKS1taHZh3IiMqoqX0YPUQdnjeTFtVo4x+Zazr7ljKrEL7gNn+/TsjPi8zWAEA
dwv5DyG9Aa15F6z3qZAA2gRGXI1u9l6IXeGWUs7J6V4u/+vDcu2xLBi4aUZivTFQl5Kvg2DRBSu8
zQBmX2GWLb8L+XRGpuvfDPqgzwkvDYILvAr9+mDSpiNpA7zNq3Sr16PAXjd6LG75Gp2LJl9W4DLy
CN3Zcr7ZwFsSlgV8F9r3ixpI8axPtKq/HSBKtT1xUlqgwZqslibplwD583Th7lFBAKSP6ubXn5XI
7n8vcDHDx2NeHiCzK7GpDdihd+u3KDgniYcZsvhA97mtI07vd+AHSzXqpBsi2/LuuaSijIpITZE3
rFj5raxqsCdtC10Gq8Lwn4NWUwB6ixClJXA66pyzJqS/oQ19VozUm4C1MYhdmZ0UTjDFFUrEtO4a
4B7+1TjN+wiwWfKvQHn4Nw4hPRC2Qqzj3qFu9ShtJLNxDWxZVgCo3GR6ZRPTIJ0YuE9rOCG3Peum
MfecbNpx6p6CIViHrGZqjg0QfgxJp2Z4bO3MAh8EHaghC6OPM66eBjMYggCKhQLCuE96M3AAI8SQ
VVzcYkKMqg4S5xyZp4Qsfq0p+F609X3b0tIXFIuAHmSQqQ2rZoJxdyUpZsM0ZDfnyKVvHOS68LSx
HShiDiXe3wLfz+el8ozVkeCGByF6PIcukzN75L1dRXL73Ty5d9K11G2hLOODSngDC/sCBUjePmes
xzI+u4MaC1DkRgrUbav3TFj7Tnf/wRfK7lZOESss08K+fsS2OZY6XJ5wFV6+tog7VDu41ntKzBFr
MPkbBHCAnDppdaEhgjs4oLF23D2e70s1U5sMmwRAO+QZVCqwm64N682+CZz0h7lwDUKMlOYq7isL
nwDQXVAkjnZ5FMqWHCOwn7OXVldF0hj8dg3VQoj+wGXSAdZGXGZa0XgS08TIQTr6brraPmk+UrJz
v0LIy1Pz60J4MhVFWG5EOxJWQJyhFYptRbR6rYg4tq0FM+Sbf2Xbj9Dn5rvg6mcVxFpzmSPM+isf
HLhpmm/zgKe/W/QdjsfossMUfsmBHu9CPZ4MS98kNBPAz0zHquXmTj+dUfUc2yKggt8cNZzgMNya
1nVzIXl39gQ6nguOx8ZLLT2q8OH6GmatKyUi9iXnHvJHAxGp6CnTaeaQWOYh3LovpkG5n1/bvFut
n/WWbDtlsRbTb7ZNScjQol0nOoVehWZ1NdMg/7ey3ljksSnN6pPuaXTzH+9p7/bDF2UWfx8uuYe8
HIToXAcX94MSTJB7kiVmqTPxTqKSapcOiiQj2HeokMM2cXmgtX+PdrecjddxZBgJcgwNV5qvwI62
MpqBFTLQBFWxp+E8QZDKe3SS98ihEblPLPSM28A6YqgRigIrjkJ4PhbPFxj7P1De+5owqHeNnb3s
qinFHECvbyWB3UqhFbz0J8ROgWslIJ+DpRl57U9EqIoYMMJ1vR22PG+bA6fRlYlZNGSejz06Jwmx
/hg6ZLN/J4prOacyOHVRR9sC7oLP9saSg03rdiznZe0BuM/sy4gIREFdUKmLN9Wl6mDk2zBthtYu
14ym1P8JpFW2I05CcVE1+nLFOnF9LZavqrevq7Of2p0/S2nItdGqQbbllRoPJxX5G6HffIY68nDE
MZP/09dWxzX6Ss7bM0W7VQGKbJZKLgMOqIXJPn5bM0yOykL/o8jUwxhFBmRqrjPLPMbz91z0Npzd
+p1mRNGfXyNue0oTtAdDDuLFJrwwd8wNXRq7n27h1A5IfGdi+YhWX0rKCtaB6W2HyZPCXp6HjVqa
UyDWsyoggAtVbXDIGg86AkRXF1aLt5pLVCAEVOIuGE9oQtvYCDmJaNPFILffIAhfwa3t7jOJnvgA
iYpeBXdm17n+3KLFusq/w6fDYYO2PJIDMfbVUix8YwKl9Vv3iFl4wRf+BRP9+daLL1+Me8svcFi6
cWCjdm959kzuBSfmaQWgng8xeBaOsgkvWxCneS/bgYbpVrWucVR7hgYzOnjqZLYwMeNh3ixi1Tax
9he45MOxYWgGU0NpLhf5cVS7fHlX4zfTNQfc9mOwk3KJyMp6u84M21Cfo014ksbEpvq0FqiKwHyr
vr6eS74tOTFRQ3jS9wOUJOVjk5COqEyIzhlbnGgCrd6Y/sAzRtyWDzEObhL45Gv9NEI7j/Yul1Hp
jkjsZ1EKp69yZCnGSjItnx1p42lup/K2nSXtpmpSpvJLAwqXqJ84P4QVFLiRWqeSjtxwLF9w97fq
U4sVMxzcKC+J2Wt4G6ayozMq7Ie8ZED28vlZAZ+h8Cc1phnQIqJ2LWtsZXZ1p/ziIGcvGDcMY+G6
FB4xYZIbSYcbalE4ZV5g4VAJw5R2LzX7NasmIztIFXBasunz/QvrYya6ofRZ0rcksP3EYLptHZOJ
+Ua7TVdPOm4M5VZtsmDeoflICDq/+SsHjATJUAeNdMUmhJOx8UM1eMZbelcvuNG4nBfvzgkrEyLM
2CANRmgiAsfTGa9m6SWyV3kehwwCpFmcPB5x7n9iXKbjVnwt4uwcFyx+zYaEtsofyRaCvIoYnE7f
EgIC2L/KGsksAL5G2i2KCjVjgUlKY8z9VXr+4U/M3RdUMo3pGQbeDHT/5Eh5T3AwaGSkpeHsqlSz
NyH0Aj+gUqATQY0Y6UDaGethvDgPdTEH8SO7mwhLmpL+7+P5yPADjj3H7Nu67M/jUTeVZUiaxU5Y
m9tpsprbOGFyoGyKz5fmx8grfueCsVAzN5cFSSI79Zeyk40f8glHJjges8Y96Z3ULR6+tmcBJN7T
eflmI+rLPtJXLQ2zpOJHJpo+GQdDeins75l+ihOVIp/tbVLGfpXU0PuPdIxpEyKcbFZhBEIqvBfF
gH5JH8euBt4ZdTYdNezGOJD9T1BwmfHjCPDz5Ym2UEP879dbZt9lmhe7rvemwY07bXsXC7TN0WTX
HHwp47OY6WTB3d4fdOf6ezKJ2qraP+rtFc/qAELTvhNgIcngxb3/Sss9GEKU3jh8sCfsyVPuP9oa
qxGoal7Tlo3IH2u/mCTkT/DgtIkNqf0YIVCr34X6XRPzxTia37Z9vlCLNQI5ta6E37eEguCVoVMW
LPi38B0zecqSSyrnPVCub+ezlyaKB9Sr+4ZfosA8cVuDH8MMQnjVAm40xvc1STfudiihlistMB6W
FE9eVNdapBowmBhQs/vavZa1rJek8pehL5DKHq0G+gMY+TD7cDmTlSAUIWLpdkXlP+MKMsXm74t1
Y9vIYOXa9GBxfQYJtFyidoDtH6SA/cR4agQl9iEmt6vq+1uI6fhgnfQlHgmY73ewD5clhAVj5Q4o
aLMuvTegmW3b7s2hRWo/JymTwf9Z0FgqrXRmWamLEWORzrsH8SYwpgkM+0eWdto3b8VHbCd1jyUu
7Fpnm/OPro47S1cBdmdAIBzJ6dfse5ybgQw/1JBFs/k6zjd2pKX57jUxYxOyWcwx6ZQuHN74lLTT
d+gfYKskTtpc5CZcDMV0PpbaKQkxckOuxMoYmCO2YniRSTHNq40ClN604kjk2uZFoJ6r8V2juS93
g1gX01pG96RrwdOY1U/J2qFy012UnAhocuNYR9Xn4Fu5p8ejleeSYVffKJfHqMpJKzwiJgogNXRu
gp3RS381JyyYSqwQN1pqfYyX8H5JzdLw6FfnodK0oRW+M0aXp6nKrGztPKKZtspXrJFKBqls2Mjz
PKSjXn0Uis4rTCRVMBsyPGSjmYykgwjSIfZUKQuE6uWLCDOWipGwPLQSXJeP5CSz/AOYqszvUXFU
PkMM8vMfIo1WZllPX375A1YxP7oAuVMmcY31VLMzEibauAxSPNgNAJwmXRDWdDwWHtAgkrQ27lMi
N4dgmxyseznO5jrLErpLKROceIdKyfVQBwL5J9kGFLzLwOH49pI8P2hhrywjJ7noOaemnNUw/juD
Efk8AzhnnhaT8ZD5OgcBSxuunLL5eZMmSi+iloR/uV2l3cSsLIlIa43zJbdyBHFFPaR+3xvGoLjH
gdf5wDF6qcCECpmcEw3s2oi6gdZRI+UFEQMXCr05mCZI46O0wTUgTmPThvQfltmUWpz4wCish43u
ixQxM9oxmXpDiyRm6mXZDQxc15hnRrbDeg/tc3rTFR1dmWpCqlJpzeeMaQr291stewFMQRXUzf2H
EGep44WNRKjyw58i9pxjZ0uxHsDzjt80/tK/mL4Q+d2TUfHD6CCTWN5TQBr8KmhWaK1ccPTtZJ5c
YJ1vzfzDybYAE3vUgvbDFF1RhuVHUwrwVjTH713MUKVKg+eT7j3Lb9TEBitpmiBKH1W7jpsG8p+X
k+AA7FkaZRXpu43UDNu1MvEcaLUmHLoUjxoEzOUay3RcpeP4ee+zjWCwMbql0nsRgg50j29l83FZ
vadlkjc+PCS4RXM9dNpOukd8kJispaEaYAS77IxSVB91gytJ2aZX7gH3TlTL7WGGESgQLvL5uIdm
6wVsQTttSs1sxtmoJP/X1v0kxefyyx6H3m6JaWHJl0VLTTnCADOTVA1Uhyhq3ffpIUO6iAPOV8/+
krwNaQTFlHb+ibktsunBjvHf3kXGsO457sZ2vxCWO3Qd/7vTHVfbFF1LczfgJnG1HMFnFR24owwa
es+5mLErfRGzGV8iLQGpO8fuBXapOwJkUHOHVk1RUM0hkG7u9WFlQQo76xauSEk1n8lmSAjHruPd
JVmOWS7sJv8AQcdb3kIz63rsJbmrRBez6Y5n8sBfrzl8tKJeiK86SkaMmZqYoKo4yM/FeYTJl93T
PTZzAeprJml2jCHD/UXjnZMG/zRl6EVzT78Bd5111uXZTw1S1oNQRnf4vxHjteYTrsqIAG7Bfb0e
Ud2JxmoHz9tRkp4xTTtqWi0MXOC2GdiGnlpaSvCn/bjKNq9L3MFxmruhIFMVFz4m6FBhjx8pGVSJ
5yU5KfIXyOiTipHD0lgKKGFMfh5xJxByZjGriPbc2fVblejMq84mkTsNpk7VJcQLaYxP+Gar9wra
3SzCgnyzpxBJ3J85yGretqzKZqUGKbdcvVaxv1nRhDj7UjCMZF7aEHEDxT5R4Yv1wiELYWmF5p7u
lQSHXUh2DBcnsmwdg8PPlzFb82O0FFaA403lZOraFr3j6aM78p6ZIi8SAEznflsaa/2wD6kYsd/2
4xCiMEXvcQilSxmbVE6oY+NK6X3f+imukr8fyXofRrwzS3YVQNHkmf7LM0rD1Sj1kwYgCumHZrmA
z6mVBHUBOtuokXnght7jd6YIazdqPv9IDPDreumSAswXUknRMPkv31wHDzECR7lUuaGbIzirebtP
EslACzt3j+o13I2vMsUuYLofAFUGed4NDL7G6fmcBalseyDEapZv9y3Fy8KX+fki6RHsoNHXBR66
GAmTA2DQBBwG7LtBGjpOTPfWZuVw8GBSll5R+RrwTwOKdskSeUJSCm3jxVfNrhYtvQbCZ9jiGlrS
/ajZyFp3GY27cccKRu7t/ZtRkLdxHzcB8rVS7ZVHQhh2LO0modfIuTIR4ASWZlnYBP8pVdpj+SzW
3ZD/srBTtRwHzbSOu/HiNpCFiSpFuzPE9A4PJx5DqGsPi+iGMMW0bKOQxa07fLrfuIoKaWQmDYUM
gSWH5giWTk2+3lDs91vitbXcM6HccD3lmVhjicUobSvfNjYHqrYVCN73ezsiXaB6djQDc1Qv6EJ6
Ey8p1yjbTKAEpEe7ltLk8OeftuzBOJ8PXWF8m3mJ1Emr1ziJy1XbsCPkfmtLGdC2B3/BS8vsyR8o
oP/ZtG5UpRHs6pJbpqM/8OlMv44gSMhLY50yTaaCkviLtS+dYSlf7Rl5kgmwryLxG8kD0watqvWD
W+j5ypopkV3kfGU1+Q+MOm0HAzmo33UsZpp7M/xPQxEzDoDB74ReWuIk0+hNW35zfR5ND28HWM7/
+sfRpKRtosRLzEeUdXpUnB+4OVoY6tIOOE4AokAq05VHFzBnc9bHVn3+qz1yzV3u+n7JF3XfsR1N
grqvBcKnStrKHlDEadxNtHYIpenurcaS0SlvK3U80a7sWkt0jovDL1njI/IZGXaPsa5nokxMKib2
0GDQShbg7TyWn0xW6PQriv9uQV5eYAKO6Oz6wuVOw0h+nEm6ugApIAGobDAPV42BGvda6Bwh6ZWW
eYW2L2K6/a3dNrKxvhvnUv+Vv+hIitFUHqmRYXgHxDimGFjHaU4BLXHi6mlQRU7liegZfwKe9zP6
9EG9TMRnXpGDIlTkTACIqr0YSYX0ZqRniFQwzG4Wv2tjpFSOWu5CHIgNLmaiIIaqUcPFaP5V9HL8
iCKus7n74BCf++7mRBXYL9m4HJK7RggYYBbS3U872Gl3uP6KDNl4mH4ToO66cch751e+79rNTn1S
fCpsbj2t+XEBJUMvMZ4KX7FLtAUTAgbK9hD+ZOyzLseC3EPzy53QA57poKBXnLGrdL4oEXmuUTem
98YVm9ZFRwB1Np6G2Mqplk6bOaOJBGcB42sfGNOMrsBv+hzogVcna0UlEaU5+YtvfaSKdmUgJHdn
NYaHY9tXOzEOvv2DUJEZlLWIurdi4zodRkg3yo4yVqEUn2vXGxC7VzJGnqQp+07BL3+ckc1Z6FlD
8kNxzIamUW3o+qvKzvE7JbbhoX3VSdjuDy10ecL/M3XJzurRgDjniJzUjOAMJsQCbrCjyE1nSAvP
V/xF2EWChuwSLNQ/xIIQgwueQAWruaR4fzr1XYwvMcgdFD7qqqX0aSo7R9V10yQCRqEDRhBxgsz9
h/lB/U7wrDkdQjwBxft610teDN71a/Ma7qNJOf5/mp2k6QNB83VE3nwXowYz2utdvNLPAJvfCGzb
mXNusGSaATxlm558Wl5qOfPpk06BHGV4BXqX0oLHmghMDEHvr/RqmSy2iaSXOW2kr+LKsBxBZWId
lzcP7GlnCgGcRfNB9782ICW46hbPHDc9AIPtk6f+cg62bgB2OaDrNGWviD7chUdcS4FpnSurir6K
wDMLT56fORiQd+bcmni44B9vZoKydNR5i/bX2dorvCEjLsL91CTb8QoF+YChzZTgxKD2UkSq0Di0
JK6QpOV9RBZTPCxQZxvQogPmwtjXhspyTnbVduiKLLtZEVF8CxsfrhDTHBTtVmpc97MYXgcn9/0Z
lYNgS7FAAWgESBvC/wSkjgxdZJ7W7VJ6caCnlI2MqpCBhQSe77q11ZmzKkUbUqrZJrFpIoMT0Oqb
/6uVYUnHogQ4vOqElPmXHAMqRp/lPahA8/wbwG4uGNcaBSkmOfkmhtZwTZv+tVG+KbRVPxzbEWnt
lec5AsFW1m+McLVX0ozdFAKHbZPOgZD4MfYJUHnp4HYqBrOT9xhs+tk1D5NAO0HFJBsnZhQ2DVGu
NHY5hJTW5RJVtCxhUZenAw3ki6gxJiA/in+uzF5c8Q3ryiLGeOfpqYxWeH92OPpV60wYGoi3VCC5
bM2MCc0gx8cYw9r1R9tr7oxRZcZKK/fesjZXG97N4fUvE9Nlybmz7FPn8Iyx4cqh4yB49EiwmyRL
fdHjgtiMZtTnm7DZvcqWpT/fgqG8LI/YB1KJfdbtd1oIdkkTVi5JkN9qXobMSM/Fe/5FUZT+jUXQ
JBmCtgqA6JMi1dzWGKkgbg0SKBmY13e9jKeV26e+JYw5pgvPYbRpLcMfq4jRLH074AMyvK9iZ0Xd
EBqf1nspOn9fXUxjrgvFKRP7TO0hCcyHkeI7UfyTPZgMsTeWWLbR1ZsLl8RyaI+PMLCYCWWXFERJ
P9lVs2ozYts5nTt9H5Pwbwwov9e9jkPQjQw1ccpi5yr5/ce2epve52JBMI9FualD7Omj5K0WHu7O
FeIpSPvcFzrnh+FrDOtORU5u2IBtYEUj01dbhZLaFEh8mSRRLphu4t7eCBOnk2CM9L+E9cQBJBr7
PyZI0NGLeVjKKcVN26NEaUGGxViLmlHT9MxOBIOJKoPov8gIQlG90UHlb76SAWRuYZ9VMJ6nbA/g
HYY0R6yDjxS6sqNsuxhgUEP4zvfG6/xuz2W4EOk5T22KzD0RkrU6Z2XqQ0o2nbeA76ro1rVt/bkh
YU/yxRvTmE3uF/hSo1D3wKw462u+ZUnTIsI5iySj2zmM2ywTyBk8K5dECOp+yWEhNb7SrvbwZYux
LqBkn47ZwjuXEaCIZwUsrEmy9NQgmT1Yl9wSZ0zY8wPvqfjwN24CDNXLezDKCKXeTxKfUqoNa2dk
fQkQkuYfggzjfogf4X2NjEQpSWb1cj4zY787Q+ZEV9uWLPIoHbaW59Njz3fMTR8iphQRrE1waiJO
z3zz8eyfuaJzxo99e1F8Wr43F5WnHn99KJpIsjwFOVJdTEE+VyAfg6wxCMBtQFN+QkSETEZyW2Up
valOIm2ltVFraU1QLbpoH5+KDIWGQiZFK9SXPkyCzTZQgKAL/JO0xDJ7s8QB4NcOJJuwxEisSMRJ
90Tj3KwaCuOq5m2XtIQSaPB6CK9knJi8J83XkUs2/wrZ+3lDKh0Z2DGmBe7/q7miIdxloJP6naO4
by5FD11QaIE9UOk6Q2R5j0+OFCQPZ81BbQUkJHQ2AYufIK9+0AWFsQZC8mLmkdVm6Yrip2wlO2IB
bhq1LpnBN+u00cyljgGpz7PWreUSNmo23gz4PSOZoEL+tAzINRdK8hH5gcPCxWmhP14LQk2NvCbg
oQdaowMlxn/CCKYpXA4jt3A97/FKHRHw//gaOFZvINLMUTi868Mw4cKzfFDfrBorAPPB743cESUN
VeOQt9CahtaZSTKfsPHLY7WKh59fB6wUM8s317wWYeFiIEcnK8ZVndmew3DjZGJdcDc6vH1qamFm
McZCdcyF1OBdvYAtculAbBfa9XLKIWr+Bs8vyvuYrgv6QJCiBYp+omu6F/luYb5/63+iTrIW9deT
ZM+wCUzjJ4MPNiK3yWGXmAb312/4gj3DkoYUQbNYaBwTWYOPiKedMerBP0suf8t1Xee9AMEAiw7/
dOSgGrCOWAyAX88f/jcbzwPppsS6OFu4BU8EXz3E8G+7d0cvE0JVOhh/8nzQ/PKK81Vmtwk+1bVf
cvYYSEZq6Kgq5XgwnkPyM7JKNqdMeoHToGKmBA+l0ND0LR7717aI46cKQAdkCr7PFohpYl4y50o0
BFQn+TUetxvWpG2mGCfQ10ugSkQ8A2+p4iCDL+xoPvWJ44fAkeHW5zNdKcFOHd5vHtzmLDFRvN1Z
U0YkfvYRuPuZN+zXvdttHs9H8yhODPuw9oaca8xG2rTTeqBASNsWfQqQZFvUl9IQ8Cb/XeZA/q27
DeNTDdx8UW3I6qnE6oXhaHlpUDeEC9HoDSJA+yiM8eluEJ7LLMdRHHRlOJLp46jjxC2A/K+dpqUq
IzWE1Pkiy3duKDt/xMUUaa/eQ83BxT2V+bj7qIuCt7d7NwDFyfUxOOaOYMXCA3yaJEe3PfCqxnQO
HBAvEGziH78w2W5NrKca4Fjz6qRYwhKmnVDZaohXYzxe6MLIElw/raIbm3NIUBQ3X3QGds2kk4p9
CffZXzjx4MeV90PEhebkqEV79uJfF5UE+jTr+HBfwr80fbKjGybM6n2fhUhe6YLQ1fjNy0Ap1Z9A
IuHrO75quMz2pO28ysa1+KbEWRxHTELtwOpr6yAkqHf6M5YBpbLehe/LL6spXeQkaUTklnpGe450
BppYGaaa1hvRok8kSMbCU8ajxojNGoRSqDM4GrgdnFvg3JYBo4zv/8okM5AJSt9Mx/BdM+wwATYd
zoa4nFSERnxxpu5fR9du0DqCnrNoild8xBKbwfR48Jmlx9V2D3qlS1OCj18I+aRaKHMhB5EstMJW
rT/H3pZtMg7hZDWe7c6QBk5l9bszuyx0yf1N9Or3bM3vcZbq60BSOiym81PSQEZrUZ0KEDnVEfDv
YMuaHI9MHRyPukLfu9mnNE3PeHRFFMRx8f4mIYEwnYOdTz7PnIXvip1MwZVwQy9jY/xdnkamieK9
Kgfk11eOZWCipSmwMBujj0jfH/WIIIzqQIDJX9rmJQU+k3oBaP+AUZr+SP9uqm3FeeALMyrPSnGG
IxhpyKTHNTpcNtoAJZBAXO9oiKJMbdHw5e7dFjwctNhFD1OX6DwQF3qOk7XX8UimHPQxVKae9AQn
KU4ZnbJ7UJdSZTBwPC+RsAD3vfQqNZ95dhKgUbRUHq+XP603APCTUU0tRRMvi3jjlWUeYbY0NVGU
gWz2yzqUysvBhgaB/XPbKeHd7KUQn+a4wQ6IKELxJU9zzqiu6H2X+ObfNPE7gL94Q1RQA56sb1Qx
yMDjSEb8U3MGg82+PQk8TmD4uCpIV1rkjBsUuxzKV8J9mJMuWGMSsZ/dAevMrvkc0LeafRGxNBud
jWMoEJyxK/NXTLwKKnd2vEFA7/ukJacH6ysIJVa+B9C4NiIHv0gP8Xwg7PrdNDeGDMGcfpkwMtUC
LW+lbT0K/gI4HiJe2nGhKUsATxPZhiSYhNaiNbOdVPZSlwFDkQb+clkmDi7bHEZ4+Dh8tk4Tb4Yi
DXdIZc0l8ctOzkBqtiANLnBgPI6ct35EOOuPxHhSGNLqFnt3Zy0LqFF+BQ2dJqQJ5K5ajXfWg7Cw
s1zTUcTgWw+cYtzQLh2/wEMPa96mhFHRyUz90BLH2JhZ72mtQSIeWeCoNfih9NPuPGUay/XGTot3
hFnfgPgdmCuYCHFkRL6ND5es5ENSyveBG8d23+hLzioRjXpk0WjB1v3BZj2gWb2EjdXlp59i+W85
flQ9RcYdUc3un0bc0QSTk/jSR0t9VgxNPgwkiLKKqzeII/6PdUJyaszpLjsI3fM0K8GUqJ2krunO
yt8I117JYBqeTbt6Y9Nzk7RT2Ui9YRQ3TtaaJQywhST1wGY9punqpF7iJerflc9I2KhVwIEy3AXK
4WlyY0KpquRuIYLvqcZKVmHZ8RfdZW3SQ3+jQO8+yh0gg4DL8dJPafXvgRiqB+3EvmZ6hVku6Wbb
yB4XLrluhrQ+UzTjsDMr57VdRASi04w3Vadea4UTliOkbZIatxpt6Zb3ziLmMxb+DZNeVSlSEv1W
rcLbeRYSpmEdgdAugMCwR/PlmTPeGo/qvpn+36bxyjubBWRKnS9oht2iGsJOzKdaOFakdD00zloN
kKhSbMQn5hz1nLD0KK98ofbWmrt3Od95EwegEIdK0PRsMsTNF2oQnk0y3Ki6ZF+c8YqDEFkd5Zof
U2r+D62+GnlzUsevIegqR1Crq/XUm9nNlmmnGHzcfJHKuUIoy9mBs+Dovd7YuzTxpEKYr1IIfTNm
KUxLDP18seSvb4phA9ckoAHpwMN1F87vTHqUk+LBhfZBPn8eVR0UFC/2ETKNRk0aQ14SiLQT1cZC
uOTBGKCffl2lpaoNFSOhTpAT2HdfEfIBwMAEooVNsszP2WYxEHN+fdNDIn2v37845ycFhOJ9hbO8
YA8RPjjc98sFt1p/Mf8SHSTvFCTL/rEWmWOH17HZ+eyjwNx8hiOg4YLG67a6ohavNyqONN+9OrS6
RnJTHNRa5LBcTRVbd8ITdB+sSZGOtdEhwI/IcKEiY1M7n1ZiQwId0UrNLDwNGWMJp/Iv7+ucH6Wa
KZhVNsr3qEpmAzYZ7haphxGR8+hBdlE9MD29lZ7rNNVZSWVNx9p7l7ZupyoA20vtpX4ft16bhHF/
NHl8kVzs851J7PfUTnhugrALGKl69bQwA9Fc0l/t66af/FczG1YFL3wnrNSryehAobBH9kADgIOu
ab2Td4ndqoRwuU31gSh89OX1VZltkw04joJsWR2CA5OmdrxT5AZ8XLpKWKGj2Dgimt2gJiyb1VyH
Ud582v9TXbbEtXLsjnLIuaDoerSc2EOdr7BNZC88Yaq6MdTq722UMO6InBQGt9hKDUrxdWN8rLY6
1S55S/7gPYNjf/1WdL280/v+cDJIvQU19aXpOGWUxVMaMd9tz6qHApXGGBJbG9Gq4isEL7Oy7QMN
TOxpCe6rcMXhIQXa1YAqxUvcf3Ti4vxO4zUZqR43a/C5AFfkjm8S7f5tEG/6DDTOwsJg3NMCLmuz
DQjepJHZytTWFSDG8iwV5A3etrRgNhuvpGFKhUw+J5F9cpoDj0YubYv/5jpbjWHHH3an8ZAuKscg
S0zKkaRprvwcRBXzf03Y/wd4wZb7BKGHQb394FhadhhxYppeawJx/CQT5GCJ+DoVJuNKxxNGpfDg
HLOum2GxnZaQ9mIHp6mOHev/7jc0bT+rN0NIipu54lWRj6tZ0ZGLPENgZHlNuNcmgK++HFMjT+DW
6kgolrTEhDHloA8lGPQpRHqcY9o0mldgpVI74082u0osdN3TfEdTL3Gy/wmwnVq9X1HSXjmPwTGe
HnpyIXjqr/pFgAWy4EDRGxzfTtFpdURzPbcxgKVHe63XAJ6lifUADDMgfIINOb/2GJYCs3nbM8rK
z1zwaTUEkpJ+tkYWJaxHxZIZv5qaunO88hAA7DDzB2+q5L1ROB3Iy7CfwlLt4PWRcoF58airwd0P
0hFaD/oXwicWBRezIwY3WFXLknpsq6t3qnapGfjR1rWVuK77rNM++765oSUwWVnBHA3owkd21X5k
rXURmW+SOrYosNydQxCNqEUp53Xphdw7RtsvkrkxwjEfhBIVnKKAt7eATZ+05HhGZNiise5juAkV
jXx4OcLd0jsEwfg7+tQCF0yV431RIHF8TdF/DA8plfskAQcRZi1Sq91n7CUwagreVo0M+udFC+rE
UCqZrh3La2lFphcszvS99kFCufDbijcRWzIwhGI2jbMWAlLg30fAWrp3TtCf7nNkX2YWcx6SSz2S
cRjJJEJnAZZ8ARRQD0Gfrf2X84HD86iFUxpNJLWzwaXzdZ2q2sHnV9ERSWtwT+v7n5o1rNtFPUG4
oMHRt8CWQvpWO60y6qsw41uL0dg2ozY101K17tdXgPFvYT2zBmzKrudUFZL/8tAa/VOOU6N6SdcO
fhJKbdJZNOpVFLPABa+SclWd47ef/upxITuL8jELWhY3MhKQCZt4p0bWllip54OCGYV82lL6CjKo
OKytYTkAv6qvoJcSdzdd4zSxNOrzkLAc709hpOEvV2AoCDwoCbZMey5i61jM1K8Ti3VvFle6acE+
AyfyrWgNa+TYXIvjSpJ9nLu/v15+IthV182NlZWSCjKY5kps5vVle3hWXOggWhmmG7wyffpWlRG4
PYTbjwsAEGm3favQQnIJjPU9PKKLhAxGcsyIDvgsKJaM+NM4AlGmSTNU/JqktAySjZMxO4ssJXem
670IGNlXXYZt7fq7nbcArdxBmZ113kFwBBjgIyi1/FGWzzyoDZ6DHH97xbWBm5Bat0q3pAA6JeSZ
HGxW8YWqO9dutEb9zQAlYfJrAjMUqAG3vMGfQSuJfuSUTJ4DolfoJtRTSkdyxZeSKFmUDBDNDpmN
1KA+TvvsPc3D4aYlhcKiIm0qCgKkYapPIQksYRlq7j5ai9GiCW4Wm1VeFd8aiVX3Rv08ZfQABuQC
KwUYqtrgSWqrbwFwXA1zYz6y95OU6iBwccJ1J9z7ZtFvuHG2A+nCTKJgyr8zCsLePyOqCDlqLFk5
chuGNdeVmC6K48U2NUiycxxMXTMfuoMHadC6QCvsW1/Im33rhzF1R3F0tiv3HxiglQGbOmbRusq1
LO0oq6765G0k68PY0qjAXpKLAHg5JT3Dk05WCG8xhRmR1stNiR7YzjLWhKr7OOcsINiZ15J6Zy5M
PpZva3CewN0VZrf/OcBmzqpE2FSV4IFmpxPwI64EH0GJV/XjTGajra4uddrUtTCY9d0DvgHreI+R
lgRDHpo4r88s+egdNI+TpuLOvR3XtkE1yNe3Nh/p3/tjjP9NKXCEWFV3TcZQZFxhm7rTG5KIzIXW
fqv2FUbWWQUf21wBP+U6an+8I+ZKdntNdTIL05rXtoAl0bhLOFTC98ZG5g1EMM7ynLsrZ1k7J0EM
WvgEV0mA1lqhB/YBob73YEG4FR6/tMLrNIGIowU7vn/r9Gh5pnSfI7mtCmy+eNO/IEv6sppZR6Ny
6VcMS5fBDp/FDJ5N1WPcvtTu5AbHbydpSkJpM0n69bp0HAwCF8v66rvSkNU2Su/On8q3UzXHbxHr
MUI+95CFk3yglbkyuBaV+5tEnulX1Quy1vIKFBph/rJNOf6w9Wx7R6Uufd87WMMrBFMwIk0QgIW+
uSyu3vgSe6u+7hxhguOpvrCPZEC6co5hiKJ0rTLOcw7g63/lZG07aGTTMpdmTwXUWQcbp5P19XKB
XYr/y7A8msVLyu+n6ytsME4dRkVmstA2KPE6FvXe2t7vRwMN+GIGE7zz4/DTBKXKPm7XnPlI+01r
WCdzuG8trzcw7TwsRTvupRBfZeN4JDKCi7Du+OmIlvQ/CGDtDUEfClCwS4sfNgHj3VBMA8FMopFK
hKZI5UId2HOIuVYwRelSeEvjAo2kzle/0mRyoty/I2vO/5cWfUVQNWAoYS3sd3fUUcdyDENnL5w3
0ViWT7XlbR6IZqUsDXAxAQlKjH+YnvDxEntYPJAaHyy32nkkthD+bc/RUZfgPYUUV0WFVyuPseQk
QHRXzA9XwhdcLKtnUCbAFupRo452r3czY1fRkq9hv3ZowYeItRzGoxvh+a3Nchpj9uDQJMxD/+xa
O3floMEzBsBXE2r7gezIwiUzVDcMGhxpSM1FizngRH5ubyTxPqBCRalSPvsyWw8PvERuDjL74jdb
LbbzsdoZVMeXscAW6Jie2+Zpbn5wiwL2JYRdLCm3xaW3JUhtAgkv+N2IrDcneOpbm2zxIxKeeKq2
2yxC2vrOScXDO0NlG0HTbhBxloiPJVNtA0Lv0gMbdb6Jc0L1QMnvcU8zfZ1wwZWXkiyPnz7JcD4m
ZUmuCX13wPJ/DKzrlKj/ycOfFziCuzznftF4+T29d+GTWQkmAa3u00QGI38x7pbv5unq1BWwQpXO
o2B9wLBBfd/M6eBAeDnDOrROQzNhFinhPfeieARq7bqvQcFbKZZxW+bMQ+lDhftweL6ZsipdNWIJ
6mFELGw2OoTYRnkUTyhJhdNg8/Qx+ktu6qvo0UUB1+TPYZIRoALiRwZDTkb4ETSkY8pqJ1aOu/td
GblKy/vfNtI4tZ5tN+z3Fa5fltBu98kxk1SNGMbwByICjsTPUEW4in0fmovd3aaDJWnJPFpdXcG2
HGSIwR5j/8211YZ4sl9PCsCtgQ+4FeE7AjtYrgPX9l0oJ7aoxb4yKKq/FyCZHq81j/LXifN7Fnin
+9PXRgN6NOUeIUMbZR69WCa9HKNmHbbl491unY83Vuo8Sk77osMzEw90wfnkwCcTwBkLashcEPt5
qqIU7GQj5OYqcemytgzcL/gtZjVjoNn3vmVr2TcZEfNSeOgIudLKEDUXIWVAgkvndYOJDp3Cesdt
7a4TBO77w3WN7ZgCTUMdFUQb44LS5NjkJxFOUDnsBxDh8REjtxPPjhej1yhYikCtvbj5E/9vn+rF
2sNfsOIpr89DB2kfVjkgilAWXQBqa0nbD+QQL4ATYoLNvBxj5pAGnTezMiQulOpUUwaqo8EwurSZ
Op5CrOwAH5mojLe2umlQbYFM4i0YnKzXb68+SSe9N6cKAdIItR87dQxAjry954oys5g5PAwZmsPI
o2EmEsPMA2Xmg1a2vJ3lvOw0F3CnLni6GTDTpvlVWysGei+j2JmxSfs2JxPTpUVJ+pMHe+CJzS3d
30ws53k2TolmSAGun7XdqZkSSrPkmxsXj0A1Yy31uX/s7QsGpL80rSKhavL8Z7JQfETtSKdgjTlF
vHUBkSUjgbsXJ8CQRFgzaCND4TtcMyMl6vxx8+33AZttRX6hxnjtfezJMME9c+Sj8KCQFhR2y1Fi
K8pVuqwuh+EIoSToUwEr1XzBg85hKdsZZgIc9Nwmpy9cLghOwsge0Jm2V0k9nyOxbIKljkiZbk40
RBAEvnS+q4zBCGMY50cGKx5ZEmyw3BjUaM3E+FOIwxPGhPfSlXxdA8GEmHfkgWQ37nopJ0joHbac
CS0CWGln/TYBfc/lCpqp3li6HwphnvqXPG3p6ZUrMAqM6Or9Vxcobew5QkVcUS3ShNK7HNbe+tgE
/dWFRJSIHrf417wZbWeZPVAymrYCPEq4XEOcbSEV5zW5nyKbjcjWeRde8cN8UIRxcWSJI2G9gK7B
JaNBqkwXUDkzKpdGClfupPGW4Feg3id516OZgQkg+V6O0pxdkIxHTTKz7JQeDmagmsyCKtIt69vN
BkZNHHNNYxX+pgjBYp+yzIheq37VRE7NEhO/YoKYc+9q0Pv+QE7z5yQO/4lybrGLK7OQeVcHZ4w+
XAHg5s/CpoNNUWGyxLJtmaFwcCX2lJD4K3vegRD2IbPBM7zeuhtNmR7wauO0PaaCkBg5HZ/JBEwY
duwvmEFX+00pU4RDLA5w1WRjekCm1JtM/KAGTLBGrJ+Lm13123lb6ki9gidPGxXawZa6hNlPfHRo
qR/CmlpVBQG3KXCfiwbu2WRga0xc/zSQPjUwpTkXSVRR9UqSAign0JLvOVsJsxPB9C8grVcq495b
sbJ99qJSZEDH6nmPRUdFM3pztXo4CEd78O6DdNWKPWoGgVF9HRMlrTVhLDEItkQZmPli/EpaKbqm
PbCtsX8D641jdBJKpyZYBnQsq8sacOruLOKq8UQ9ipKVtx9FyTNmdsyohccVdc5SChXfZQ7kCeQj
UUWO69pshwkzK4MMVR7/gJem6/0X+E4SANJ0C3bPJiC6YVzjutkZ/GVocFekWC2bsRAfI6HDIXe9
p7E1Ck6pKTIZG8TTG+yAvmAf0GDRvMVgdKpG+7i/nnqujFbqM+ADLARtiifTM1+aaPFgNFG9T/iT
+MrZgRc2T50rSEZEZyCqvurWJNVh3i5mF5OMJqxrFnxRDlSs/vUeAWQRpGrUn4fMm8zoSjQtq2du
p/lSrbUw0sR24Req/FT3nbjek0txUwugPGAWnjz54bYEWJ7b9JVBC+5JHrBjlTCt+7hzHvMPjLLU
PsyCG92s1WBqfMI7xSHoe/Y9n5ijLkljpeNhDn2KDQ13AO6NRDJoo+i6ZklEJus1/o5X8yU2kS1N
nypsaCP2NoTJ1kgEFqRUo+i7wBNRGrDIViD0tmzzptTHRHCuVXYh0HgWT4BpiAOEq7MEMfTesayO
62uNJ1nIkWwzOhj3fAGwL6fM8KHoeUvsquxMv7pRo//qDDG9/OjdDRSrbSAVM5UWhZsr6lLvqC5w
VW4VAMc+hWgEaPl//OeOcZGFy/BijAEYhOEjWVg2sA35NDxR0NxL05FgE+NRarhy5Vb3wY4HSpV6
FTJ+k0GlqcFoORGuDSNmsBVT3LrQSpq3Hrq2xcBGrf4iyheHBscD3NFYdgsleZYk0DR3Bngfwu15
lPT1j+qtffl2PeTGCYxL0TB38MGQnFZpxZUKsNCTqNJl2ZrspSPPNPKxIXMtPpW6IXppKgcjc8TJ
ILC3KTfDJwXKF3O4chOiQDK+jKYckMQlrDgJD6l3R+oQOGzoMXlFKksChb8ZHLYta5cN9f4kyHLl
oaNgPlebrk8N9/5y++S69sjqhFl+ipdgb1EC3YLXFOZgnTCzBr7jRaHHl5C9/ZTAfopp1xdGTRgt
KpnezK7Oqx0QvixHW8+8SRX16EWegswSaj5HxM/hqssNwtXfNmyfb2DhS0ZXEIuDJbDC5EASbAZU
3reFGpXFZ8+aha+X5nhM670mgk0tPKdE0yiOXIv5A7rUNrM4AuU6wEyPT34m+4kRKBSMz42PxFwu
tT1EAHJPdIJ1vFmSqtg3FnrcoauGsr3dAnMIbfCooCkzq6ZRosmLhtzHhio/2EHM/wYdPPKVSDvh
7UixmB56w2TWhoD2Qq6+5US9zbMbgx2VchCaMPrLWx73HX+Sx8MTKAIOw9fOO8y0JCAPFsrIkRm9
zWiYUz9lL6+DFgZuJANn15n5uKv4tUeVIZO3k763u35f2/rK3is0jSXzL6q85arL37fz88sJciFl
+hBMzns0qbxO6bLfONf2YhoX3e9fPjKcnjAFL+sYsAKtTiYsyKFbfl6/IZ6OSZnR3dVVgH6R8RwF
IoyB2rmUqK3ndlTG2CPJSCatQ+S5JmULT0a0eK1LQLkDv/ReueQ+E8lfhynnCZ+h2ERYFTLi1ehb
UUMM1h69aLZUIseC0EJGD3zbDX/1DpuzPJvet0wisPFjBKONwa7UJ7tDtSEj7VIu0U4ubuPgNu61
BNx5Bhgiu74Y/F4jmcykBAMMQPgJFxf+tQ7KqubMKmxHezcLiqWsmC5xSlwJQtJO/6GOPSnqMd6h
XerY3WUH8LThiq5wAj2AvMcgdMaI4ZaLVdwYIbEficKkL0TPGnK3HfpxAfjluzQK3PbjgzvFMeeP
N85S9GPdVWXspKYha5/p2Hg2dh3qy20A0fDONlAYdal6lHTrQnuDI1u1gddPYL5otKzPCox6/vLS
lp5J3k+N6p5leqhIB5nfCVBwyDHDunQ8zkS/C2/P242F/UJE+XG6u2gG67uvo+tfj17nStDeHJfT
HWUcBQfGAMUqHoRFS42EKjtVtQGzQyJxZ8x+PMcSNd6W4asOiE/SoGieNh6PNheHSnF0TSKV8+kX
0rrtaXIGf48E01+XRG8hfpKc9BuCL9YrCLeZKf85P1AeHkRRnAOBPom+vX1hRfsXAnsyjFypuhYq
oe0VRZpcBN4OxekBPKR5HQAE5dsoxwU4DjEd8nJcyTK8I1r6Osgv0dIypPEfrRCIuadXLiS9TOIf
iMtDDnfAvWo9CYBoyxCibACX0E1QLnPFsaVdMZSCILVs27x+NoAez/rQquQIKi7Mmc6YUL6x/34y
Rg1HsJjsxg8J6CSZUui2ALpaM/u+LBfYLkEVIcnq38gHU8fnBFhzRHbXpGTuPK1eqAzVuTe+BdTF
wtwEL7VbxHcx5fxTe5WvZh5NyLcMgU8QHjW3+ogFpwrR9apnrHTuPTRvytGt9m1LIRvYoy7+8/Ru
FIwCOQj/qVFz0ktkcRrb/2g4RavAzG9oBenGVsbaxH6G/sitg99PfhAdA5nLTe7v0DfgUf7p+wHi
QtExLDaQws76fHxfgUu8E394CkmVLqpOCrm8LU81JfLP5hmKc12OWX5RyUrGm6DCjkXuaUv4Nsp7
GcUkO8C27IaX6SM0qTsjtHFtv3Esrn8hzT0McGtn6aD0IbNfv9hwbgX/56dWzMW8GftWkigYatnn
kvonX0DvRgg5CRSERwEIc+6KdxRiWM69vuPG1l2Oz6XwauzJ4q9cQwQBF4xSI4oufGvDcW04/dEF
e+/EgsPQmaBJxbfsnOyLCAf05/RFQqsaox+JBRxWSLVrWSyXzaANifUiPDg0Lc5HXPKd9YQqr1/k
E7XgDb3HaeLze7u5AKS8vXyUTt9MIiajDUPfYu+eM5l2C3GFc/ngcz4u4MqUNktXt92/4ZI2GVlp
zNogavjekade9OiCvNtF940ZuANp2Nckb3M3UAOWo/bYwn/dZbGk/4vACVLVPpX42BvhhLMT9osN
ir5YWzRPaPq4tmknWmFRfj42C7t0/AyycBdxNFgOf0aLZyl//IQVs74i+JPQV/GTHaek2ISWee0/
QL4PKp+NXx8gPO8ZyefaXLBW3UQmZs6syEg24Qv+Ka7LUf/3VqDhDSDnBa1543aL740trxieGjnd
m7O9V13TR8Y02Dtaukpu0jNGoH9XwoHbyHUSMFOL6O+rvidf461wkbiBN8FCh9OGbg8Oy2R9hctV
yt8FKsAdu80sOf54IcgO6L1sQLusNUzNKb23WHfGjB64C1kyiWrtT4x7nd26z9j9k8OW+LrO160g
DOxd9o41EQY73E1GTpwoigY3z4MXhD/UFrZ/cBggIJV6qqXApuPE3pW7meso8hpmtV0d+N5ifvNP
XKzYEL8rJAA1tmuj36PiQKA8RzUEuuMD/TV235lE1OyoY9hr11LlQitJXk7jcA1NWEMMD1G6Pf8p
CCHV19dwQPRoXtDo4b+DlsEYM8bPA/4Rp5JFnx+MQIRP8/1I539M9P+7jJRRCIxlFn/td1rgsC/1
iVBfYjLnREeqe/+UL6vxrSdzhnWcKNZlq/sFh3sOAFCWyAID3dnaNvxUDDf9ZO2aUluZLIDel6ER
whpKmmPAFh4ijQ7dj7VLDHO+DKccvCUsWjndw8GFmIEl86I/Tj2Qxu+L5+2FKkPZeY9yZgeauGIx
ZsZ+MaaqK3FUMnE+E2gwQuSNJQjJRJ8NUfDHpNFAYX34pjw46MSDOZVRSFf8K5/dA6ngDWgkF4e7
TyPZEoRjVEiUu3fqv0uVHwt11n1ZkeazVyK0wRrwLMW4qovvBkoRyl0GRs2jbafCeas1+9r+PEcQ
y89zPwWfEDz1eTEKqUMGPH/CbUkjORAw2C0Iv1Uv7QyXWu84nE/EG0clImiylxbL9k8B3YmddvJ4
pxDtGBRik/r7EVEWP1Fr9vyHhSN8e+9uYCdWMOfXvswdEZxqAXq2LHtxFLyvVaN8tlP2p+VsUtZJ
/9TD/7HuRMWz5ENW2RN9yV0dBeBGMQRzVzQ+sSmbALwUWAmwO1lKykBgzr4f0AzbYrElKgf9oxMi
jK0sDwFSm5Pvpi++kVOArzaZcqyuQWlNcs4KwpBZFR4x4rKMu9OoFHpSaiy4aMA39Sy92thV3DJL
Psoc52w9OUTIvEEps3B8l3y2befNuPnuy8t9c3AbLR45t2Qyw9JggBfnHN3VuGoo5Q5MC3Ji44Pw
B7dFGTJTS5BMfidiQgnvojisi77U4ezF7a/akv8ACj4l60ohS250n9m8EBonppAA2sWFDgFCEMM0
16+LvG15g4k9HG+VedN4WgOyw5iHZekB8zIYkLFSihprWtwNPkXZysfqsrABaWqW8YBmk26Q9ouH
oAAVJiU1shcM9t0rXaUFM1LKdNFWQ/qlETV91dQAviio4KihHzzruc3o8/OwBWt4pZiJ+OPFq5pt
E+OWT1kpZL537Sgs/6QMOHj5Y5rM/sM71IX1HaXzBKzcfBTZ5ULYFJ2ND0dxS/0DKnM2BXMzq/lZ
E74iEau7CBKDvSIUMPYyuVEWnnlVW5/0kB02IUt113m8SkBtTO6hF6Ez1IUBTC+E9yz+n9C7XBuo
2ciyezD1C8PWN+sZ72gVnm83ubKuegtyWRavkmq87htmq5TF4f+mWssXyit33ElbHU9dQQBs3g1l
XW7ELjzl8Gf3Oshq3g+qQT2vSQbnVK+F+a3htawxRlEgaHZioLnx05vjAXATbXMPysu0LNxa6cXz
zg/1AT2r2h6fafL104PCxnYuPwUogJKqiOrE0ABnEE7xzEyFhRIX/M0naSMA73Vv5NSR+N60rrBX
z3AaI2W2O6soqazqtfomdBbAOaNDE6PwbIp/gWNqjcSF5hlvNmLYGDvz1ABW4aW+SY0qleJjSUcZ
LKy1RR0sEjPuerQ2Y8Z/TzPCd15lCLQA2rTT43Tj/3U0dNeFk+XJQb5VDiV8qPhAkWV3vowzxsc4
Aw6hqLNVu/XFdnNJ4lUTNiuNVlRfj+iaW+HOmzXzSl7REniMh3uGs56aiLVy3bt82JvHl6EsY8qj
mKDuhP4pF5Isrs6Z31hJ8cwIrHOk1dNwKRABt6ZD9FsiKJPRSjTOXz0RhfhCE8XtMJDzZ8E15ynz
2pq1qhUdAhxoRfj14KLxedUPtzhmfC+e/qG/TH7wGQkGmV4fMyCK7YGv9KZXvWueMwsFd6MaCLmn
Zxy6TuZRKAo+NfmoRIHIiThlwDMQ/RB84ELg32kN65QFJaaW2sNbiWnMcN0j0MTgeaAL6jA/vGXo
etfnHngswD/jcID7xP6IEpV/PN7wWyUaTAn4z422YJOf0ZMY2M0wBtPiSEoEezUHuTDgvKgysEvn
KmU+DzcJNOCZJWK9ILWxNS8WNVtq++nYGEvo1Zj7y36Qxu3cdeGafKK0y4MLkzxYo2nJhvebg0Z+
EFqEKWeQt7OIbe7iQa/B1ik1BEDIm1VHJaytWJGLEFMLfJRg+bVI353/3PwNOqihosLK1KEJQcNY
dsqPjdMWKNTnRceShsVXCs90K1aQbcPewwos0ye8o2TiT/Y0/vn1bDJ9ikmvsiyZLoNiJXzXc+H/
zF0/rcZifOlOPymVHMBwR0UM7MOyjeHIzm6SWuKPnF2siW//5oZkY2plYS8qME5aRXY7YXbs5nFo
MDPB9AMKPR7L6w27b0iK3c/wtnPZ1LaMQjMv8aYepiPjRR+2nkoH+98k3fGwivE2l80XqbhhUJUt
ihzCD4CUnwvpvpPe5rhzamMrrOYocs1ZyJJtVq48ZcvsR3mwGSNY4fJL26Broa/Jg/xYu9n+q2Vh
s7cOtyire52/G5UKgBwi9QUYRYulVTYTdhgl1BI9J9Z4cPS6ymD7mNYcSzQX4Do5yIyhhU8bj3g4
feMU265Oa0x+kqDwe2YxDScwcNYzZtzIw16MORyUBicN76cpPOvSoKBa36qjYFTxFetzqaS4hqhB
shAxF9nuQGmL19VpUe5PrbCf6UY4RVNaE3S9Kb9jHQ+UwNMQHYSojYkhw0W0sYVs68nZv4141Ppc
Edgmt6STnMbcrE8c36pn3hkKmd0Pa4EO1vAF37A0WC0B7LGI5eTCLGgR4cAON0FKfzwLOaewjeZC
I8r5AUYZGWK76669ybAsXDhd5olMmy8Gouk8MYHjeMo6U3GtZ2np8qXUkWOcyjSeJTTXrLw25ZTb
5Aj7hRY8C1mfYjgaS6OBZjpXK0q06C0w32u+Ss7ZjQDqf+eDpdafNnssNsJQ3a3g4LgYk2bEtfCD
HuZyFiGtxMWvyIsw60QJKi1B28JT3XiTvmiaowOw1opOSU6wTwudDqpW6NPtFXynMF6x1dH/tJnt
NkVvXDG5otEAlwkipg+PL9Mia36MrzH7pJd1OZjz8X70Vycl2/Uuh/eE0Hb3btgp9n+GKynMqDDG
euh4K4ZBg80LGmx7Wq/pcUlcGdMiPMYdcmEaji/KS5nMOCCMnnfE9SDjUwS1fftjUXWEOLwp7Ory
yU7riPlh6EaKgini48/PawRd4rO7zWQ+BpU4LLI0xtT0Gw63IygRnuKQfFQ7cshBHTVymj+Oh25Y
cjWg5ISimab3/Xhj/wR4MhhhqZkoNjXzNG1Dn3QFHZuSFoqRJGl+BpBkywrec1l//Kd9sRQ5UteH
x0cETlnRrkvPcH6PlAQgnQERTlfq3cKRkTBrYAet5khs188SctafL+/xcioFy1WWGJ2ixAqHtnbl
gVZ9uP3srT1VXNWxE+0mcAyKhtzlWUfxiivRa1NXyZb3oKBu/7qXxYKkWRl5bWSG3n9UevIBOCb7
6N454d67LE6cS/3f0uH4VOEbSvfN7BH8U6Rqf8P22PNJ4KG9aVUKtLFO3WwxiSD6tiAXLCQlOxnT
XAj7WGHSYT7jBwMJreQuBn2/UNXeORu3ms36ynSRuM+DD4IGNvzuPEalMNiJQ325jy/ou/qTqT7N
yudvgAaCD310HQ4xBPpymAu2PK7qqYHwlRlIE2iQUnAvFg628UhTDkHbZaQFrCxrRPIH0jedqh0r
3WeVBQL5+DQZ5Hdw8XIWhD+zG7ybl2WBjJQPnML1f+LxUXe3y1hPcbEm8eWS9qTXYBk735fBcUV/
gtGd6i0zj5i0AxByoFRc5lkiRPK8sGFkTpWbbckW9HJ0QQKOtP5VF+ttadwGMyKf5KZCrJUnCZOh
OGbtZnG1m6lzBc9I4II3uw+02oO6WQBNAHdTDqnvpQIVMKtpicmdNCpbFWZ2iLbnga7+Gvl2Am1/
MjunltToZzkp/05BbOViyetsHb6t6cw9bWj7rA5YkPjZ0Tczc2wgXqIeYSiu+CNhJg2bNjSWs7+D
LMU2a/1Em8SQZi+V0uT5XQfzE0qe/0a6m3upxVzluuY9RJcPmw1Km8pt2J9hS+ptJtH2vwvdOAba
PoNK1Xqlbnq+qYIdStKLBWS+qHVpB+1e4d0Zfg0JYhgKYFlRIsard5yT3qLuU92MqU9tukkJBw4g
Kk0Q5DAD9ySYtb9I4PBJh/AmRW7dZzmm7gtwdZkEJQp5GSAm+Gze8YzLF/yhw4sACS3gzHuUg8Qn
yYzenkmn0ql1F4sMExtfhfVripKpvG8XHyMXLAbp32o34EVb+xEWDKRSFa26fhcypFhCOh4S5X0/
W326Df7wRN+57hYV58wgRfaZrhECyojatBSRzkJeLZzTzXwRF1TeMHu53Hq/M8tfbD8DGFXA3d8e
PR0ndKxrC6qtHlJ8Y1BEZq35VXiSZvFvrygaMG+/1k8+oaW6oecj5pFltRyVGfkfo/NSIqWGmcR6
SOYqS2bddC+Zaezfzh8I1ownKEs/SMZJMiEom9BOgJ6H2iKBHMx6liAd/soHDT7f8WfciICUCd2I
yG6xR7dj+JqxIkm2cRXtXBI8Btix7Wk/yhcG9YpeSQHXEGuozDGWSEKRUY4sYLK4uuGlQlZjddnq
fNT/6JHUAKf63swBhkgMR3xCYlO4hmc3IQ10oW9b+JkGkJkJHw8AC6YKHcLWH5i8K55Mfh0att8m
5puvUMyjGg2S+j7ahjWhB28eTV6weDx+acveNx7XqhQA/fy1fI0MoCipByMDGuBrXpBK9QvrVRiE
0oUqxrNZyHQPDlKrjahGdP3ERdhWJU2YDPA0UnYuteiOccXYaOYuCeGh1cYGbBaOcXdGE+YKyIZ6
ZugScV95kpk/WbUne/eOBSbM+5o8N+ePvSueZ+CZWYHX4ORA/lHI68P553KoQ51YLIT9EneWEFwe
b0p2mXNhhBRcnHkbpaH3UGZXkV+bLP9QlhqXMJ/FVV1/FX7uclSAb5cqkpk0JsDV9aNvZTqa3MxI
YpFiCVnRqOkXT7Seeew0TuNZe0/Q9TPZ4sK3GGQ+ZqbS8AOa4/kAPJ9hQEJ89MHFUJJlXjHyFR3I
zl/PU8ZxK4MS31DZnZGSgaozQp4mQYb7xajmVEJArMuOSrwVHiuaAIXyzJHMQwvaQN+LYVGA3XvD
lp+qqzB8yAyKWQCoy7ewhB1LFiVvu7U/eACIzAhZesBbCV2pSnnUPyS55tOgfj8KOX8zWxWzM3z6
WITFt/HfMSTAdprXQRcQZjRR8v1oc9XWHrnv1HGQ+CAo+FGkZak2/cYPzzkLYZ/4zXVfkNFvhTSa
1NWpy5AI3QQU6VXWdOlY+Y9JuUQVl02BQPZquX8ziiSoqZ5mACSOKtOgK2fVNRe3aV6vhnUR1MtO
xIO4TeCN+UEW1O03chCSQYv+a5d0wk0PpOjCs4SA6DwmQsHcIcpdO4eHZDNPlu+3YWgZFLqVRoyq
fKmOzWr2Ie45fjW1ge152ecYQiZn1PLDyUVNlatGu6JPK94DPubwB+NwcMos4DItxzIVZAPMii97
VQod/odyhDafpEdydqMC2csMJ0PgfP5jeiA+//AeqbSe6scrfidBW8RLZa778wKj1IWHynXZJkKJ
28r6igfE1j8pcd4jQBpWOU8IVU6LI72CufYk7wEgtGAC1JzswlAHD06HjKKa1r4Xeyc7K9atf78n
PqepctxMAdimnx39WFNhvWlMYt3zYVOuUoTzllqxbfylWE18JSvP6ac6m6N54PH3QejerO1TQCUV
4xd4I5LqLgZvTijDdY1A9tn85lQrlzJ4dfk+XVWJ9SxMOR/CsiyQSkRRrOveFPpnOXQRyKebHew8
IvdLo1WoUwS2vHebtPKYtfdFmh+ndjIuvZnth2UXpTnB1tedqH+OhSoGumy0VwZQWSCuQHtVe3eX
0mJ28Yxu8P9oZr7IdZxH/CzNK24w7PCIg0uolufVHOe3ljqKVEGZKQAvW7ZPhn7B002FAOx5GzOe
pwLt5KMq5D3y3lzOikhxMwdqq0Z4kd4898ShcmQ8cauojKoeu7/hPEZ/UTBn6dEwPYDumXUvNl56
wku2ERcNIakV14IKRTlXsM9WzGiKhgebtPiKPJbzur9RZO76fedfsBMQgpFXH5Tei4U3vvMMN59w
3XKK2w0uUMCPStda+QrZ0fRRA6Yk0aP7pUhTzwY/XAZq5uogOwPYppdGlc+eYYseFB+svvhonlTU
lFTHPABM2SyxTnBF5Md7JPdm9iqEbMx76y4OZNKrvwtE/sUVu+cemiMA3O+ax1HxfzeadG0Lax5Z
0r+RmqNtPrhwNSxgchL3f6dDoPcncDWo28ssoDO8c5M16k/f+r2/YlWhjmhRrw7HZduFtc9e2gZf
rtPPiPkj0oOisjzJLpzFPOsYGbhGm7ljh4EyQt222zJ2Vxj5oDdi0FVN20KX1xdMxwGVANQMZcle
i719b8g1txMkfyL7nEg+eLwEzRKsmnt7wg/RkI55LsgsTURSBe9LyvUlq4OXgy2inWOsK1WryoP0
JAC27wL9HUumXHJF+c0oBsrkvDF4Us4DkENK38DL10GvvHzE0sOC++soriV5py2S6DGP7O9RbVWy
nVH99Qw0wdEvtVfAls1OIRYscN7ymdGAFU8fTRDL9+fxyM+RubGuR5T1MdBdM4Arn5f4gunTBiQ8
JUbVauC3Iv22wHIrSR95/q7c+GeMvJCqUD/XRNWNcuTBn/eCyzJ8i8z1M5OKiFvMQE89m5+h+2+o
B9KAiGf3stKHfPMLl6YzLMhOnH/BdJhA1CM9mMkXExsFfWCsm/U2uvNUBySRI6NtPtZiol4ob4JP
qIG0DZI0EaJpzB+IAfxi2OLQjkDA3eRwNVxUJxQCm2jYB8luh1CQki+t7b78C5ZROMygthCsnSeR
jijtif8gPVCa/cqIyyg0L53aD5Ei/7I1dvCAX01x/jfqFLtGArPTv5trMVhYWxQnMTf8CT7l/f49
YmLX9AZxPO/vMOPeNc1AfvGAKm3/JjmH/AkI+idasqQAh5rr2UfoQpcjXLytEwV1HZDbv5P7ygIx
j4mGUkvetphlxHC3w5OxPhHKLWknReHYR/JzOfvmqPcNqsmoDX5SoikwhVSgtmMbNLp+emYIfdyo
Joi6g7cD2tsCj954mZjWYdbdMOpsWJIDI/15zl8cmJlZo+9UqXW1ogkuuPrezzLRW7mnLfsfDxPa
vczhbtm+4C6kqEUdhoh2HR3flye/HqbAt5Gt5dv4EwcEkasOaiTz2zc1zLXOvUW8ATln63ZeySWf
JbyOI/dKstqZkXObdzymaVwa2zl4hkY4Ddsyq2JEjADabh7wSENsPf+4ARadeAfK6sHyaDFZ4Xz3
w2HEMXR4ZmXEZWkkouigSwHOB/2MOceCOkfGQwwYXudU4yufe5iEXWNAVDhWgFcnmSKlx+o0pXbf
eEPG6wxqQzPL/uGL1wjacmUFUydkGuyK/xMM1rydPD9AlIlKO/KOtGsqtMAo0h9wXMiuBoB5h2n5
EZvAbejkeJ54P3HXqFRRd8CagKW4SIpMJdVRN9yp2FLzV4XBZ+mp7kkulNUhHnzsUSA+HZNskNqi
kL641Jnp1vVNj1Sy5MM+F1uZ1MSwmupjjEfxgkDLK4LBNZxaE911oVu1dT6Wgx7bj5wFZZHNklHe
X4tA4o2Yd5BrRXEWlS+UL5dv39JwbY5039+zSF6On8307bo3/47nJcNzHYMRCi0Odc+Tp4GTVuTw
r6J4c1e6wZuu5e1vxbHavyNVwMP0XjpaejGuqLjwGodJY3SeI3fGI4GUdVKOLosI5J1RJvtyCbuS
u9tn06wPxQJc5QoJiUHI/Nxnzb/nukG2ZZRv5Rc5URJ1ZREU1HiL8l3k3s/6NGtSk04MAv3m+BUA
8K2IzQOQpGGcNeArrELGpA2irnG+W+n/8ujMl76RojccAemjYnxaQZ6jm0osFY93dduDxeBbeFaX
751tu8gUi9uCgjR/i3usblAozN9qmGLKUikmvdOFc5+yHHxmi0mLExg1Rj9yRKFqHxNkN+PadOrT
9xfLJYyAFkHoapDcFkZJZkgLeDU3+8opCWYKJ2dsP6ZsF52rGCUUTmSaMGCnTINWOBIQPjsoeT3f
HLCRxb+xetYqCH8Kr286B5MkbfYs1wbKK3I3mjb/a6lX94rtAeR6NCiyzBr9Q7XWtZ94J01pNw6y
6M1E5Dy/hOezLUEItCKkmhDTrtfnX+YJrWVrPgxf+HBgDfLWvJJJG/poCn1LPysrqwNM6BQSQjk0
7QhR5hJH1CMECj+JCDf7RcFkNdNASxdiR6pnWXtPpRKUMlJel40WhDoxQyudp1Z3fvx9wifizn+B
kdPrq1C1ujLYsA3nLob1z7Urap0+zAEHf+qzTLbLDPRpE3g+1DgPLvxlFXzyHERvAqLneLUVMMTB
XJ04/oWcM2+ELKAjQLO0+30x7eBmkMo+hmVGAQcgwxHPfe7OSviwq5VgnxBXDgAjquTdPNyjlY5P
oaOTutFn9A/Qvk/u/9c41r3Z5boZppi8GnT/0erC/1fbvmYoQcMJlRDfsqV+yl5n6MDJvzP0zbwO
pGCgCWuVrCS/3Id6O/Gkjg0UyrxhmHKyGZAYwb3NgUByMR0BUdHi6PpZfzwA8Sy1GWtrk0yF3cl1
ugzh5jPU3b3OqOqcJTp4cYTKfV/weJoYYVRdsK3PA50uusmtG3ViMah/iDmkQSWlM5KoxlteFd85
04PP/mneMAk2+X6RyJ0H2jUleRAxJKRpAmFw3fW4x5sbN8sAPlK0IqO6VXP2lsRJVbiR5S31/0cz
Fhkm6wxorcdCbEJ/ieXVD2SHjh7Z7FRsZD8F2Vaho8LrRvH6BouzkGtV+Daa20apeaQ/wbx66/5h
Ok6P3Y2PYmbRAIXu0XkJo5Xp7ZqTyrSCcnpmX+XrUs4MRdrJyWvg9D/zqWKNaV0fZwVVbjeOZVwI
Waf+QENYsaZi6jfr1+xOTJjjXseyezJfxtfLuHH6rD1EuwNyHOaafWfKJLbA9Y8R4Bhk22El0Bvv
dWVtJMUbwbYUfQSPuVUAoY8dvO4g+jUitDMFqqXewSkekmvIWTyJitax7q8ZYnWgYiIxon8NcztO
UmaSCvlmV5aJ+TpHONnzjMrk65RL/dycLraPpSwwuGucQvwdFGmwnj8vEdGWVPJwoR4TMvg09GwG
2PuK4XaGKOkWJmuMnjs50W5JC6xHV0IkYRnBsBw+3Ko3m+024wyJTCgAzFI9HFPaQ4Ef6XHlKNED
96GeBpW5asnoTSj8bS/Mj7oKPeUypazp3elNbpuFra/lvgRb8sARAqJ3ebtuWCC90a2mjsZYp7J3
kzm1DMG0SYitaeFLBTFowvcouYg++LOEhxD0o+jmDrwwCBY3QJ6ogVm0vj/7v5GHLRDgyVWl4Xir
4PdSF0kYSyL8OighAbooOpTJhECNFf9NnmlWRFmCbtm+o9/DO5KevGHWc302yzzCNagNUa2Wfap/
AlH5yvUgWtXQhsyKh6IT/KGHfBDBZKyMPYaZdHI4sAtae8sr6kkxQyy29YPI+sNZ9Zh3IczxdmUo
8uYTzwpnxKGTr2LzCcOINbxmseq70Os5bYWoideA0V2TiVuDEBmeRdn+vfGzuWWYb8OFb0iNJLDE
LCFsR5++6KDKWK/On7zJmSfdjvFuf3zwwnwQag9YTcBLcxaU4aBwpxxP8dhEYHCQI+zXl3brJYgf
jNSZYK7Mvzy44prH05UgwEZ215sEAG/zJxGFjYcwh7uqXHjCXimFQPOh9YZz+tct497pTc7JtcN5
jvLBpXYiuBp02R2w9q+dscUIwoPvob09JV2DbqObMZ25X2uOYLgXwfUjj3IIpE9JgB5B5ptgiE8j
wTOdqVCZuSAe+/vRW7+aXJYFUr5tvFz77YHKZSbILlysP6fOMYBpOAGmzjIsPkqPqmF1WcPAjpwk
6UXAsWE4BxCz3hgakMjcAgw6ssAFI4D0timYSOsymE6HTTJ//iZ0xldXcLqL8vhk+8QXNPRWaAly
i/8N0Dr0w9NHj6sIdFEYkuxLjBKNCMvjgu/8H+tA866hImzv9EM9ah/JiPeLOdogMXGBZAJbSwIF
s+AxukYi2qMLEunVmkpSRLIqcDOt2ArK1WGraUhW0hh3gsuR8L1/C4D2z/MdH/vRcwOeZZs9uLnf
jRGtpaHTTSBwfozuXfeBBWAIww7ElQzeamdN0m57P27pQGQhb9tbF5IBdq5VlBS6UV1y61TNdw1s
YaWRXZBPkuxI8X0/dq/JWoSSK+lA7xIW8kMsQnbbF5k49W4XQuCZ8ZYhyGQRYqgkFkIE5723wj+I
F4BOqGh+RnUSFeFPqN/+Fsd7ePPqzr3RIqfKwrZ8HWipAPnHxwZUh87kSwieu0UKgYM+/AcA3moV
53zT0dlcWXKEZM1zWIi27ikMKIILYgFZ9r++Z4P41lhgoxqi4ZlURuIrcgiWKsCAPO4avK9C0uQD
NiYwS0NdG/P0qVTFox674V3DQVEk6vLICkyPmAg1jbHOE+G5JjHG3TWQjhsTqCfX/0nKROWhutBl
sMEcFlSkms60h0D+M1aVNxf2+MWzaLC0BTyxXRr7EvvvMD6cpNjx4+bz0F2jeZ6AyWHdQzH0jL2I
VZ4lJqX8Yg2+55W4n8gHnt8rzGt6ck/BgeimnRC83rQmiHU0OUbet6USkAbHnPf2GeaoBqoptXOV
krkY09rcYjDZ7011htqVoWORbV2zMJM/wPctyCJMmmtbywPFwYJPc+Y5YIkoXhA44UVsh24YTsuC
5rwdpXNTzaA22BBqYIQuyIcWYJxNBY8pfss2YkZR3LPXFXqumKonqlBcbJGMI2eAp3wkD517Dozw
NEXq1xbfZSXla1up4gxXURJxaWuff1ccS3DJzvXdojI2lwnMQWmqQQ7fr7hM64T0GERBdC/hr4LW
GxvJ2G9f54/Uv0Lhj/axqi9j6LVkIIzGmQv4+mNBHussDOHQwWFnCQm7tI6bwj0JJN1NB7st/Be6
GYCpJP1p2iamoraQa9Y945TVbWZpm+DA2LyIC7Gb2Dn9zKzlP21O96YTotNsQV8Hc6nvo8PwRbdp
5V6Qr7qkJUJC+yepNCFnVo/UCM5t5HZzEX2BIYowS7jRmT0YzVMDIo2JJKEaH4TENE6vLuxGbIEo
AyuPldi3xHDTa2hlQbsod/4wKarkI3DWns/ABvSBaQkx53K6Q/saAF449mE7++BXDE8SdfTOL5Ws
o4OP+E670jyLZSupDOxmtwdYecQeF7M1RBWvZYzol8Ni5JqS3yRtk7AD58C93m5s6askgamfm4OW
QuuWxClZPK2TEM5vEA51gykc9NUrtjc7hzBlhKnGAst/bMBTI1PwKEDKfLOVJW8fmB1g7fOd8KP4
gWWUu4Ht3tr6fhdFeOK2sJFjYZa2j/f18xPU2QZmf9JGV2+NfdD4SI8V8ckC8FCkCxQiAVUVRt57
H7xQL9NUoVK7XvjIBLY4sMJavJ/V+r9j54+zWvMBk4PnHGL8/0KegtZyevf3xBHiXpiaWKM3Sttu
wLRSvv+xz79zc5JUVWzxPLwWOTrO96GXk3lBDs/IcHOc7ZcnkuEkpFp+BUKzZ1GrtYa6YQ8bx1so
Xt7KSZjaQS3yWYpxBSMa39idepj8sUe5UU8QRYtc2ctwtqz+Eagb0L/pMSSB1BJvBxZGSe/5zhil
JrrHuN7eBfJ28GWEAqpgFnrvqcHzZreVLjpKO29QFP4E+FuJPnvqpP0F4MnIbdswvhELnsGd0VUf
jnLoC9zp/z7SP7/l4gYHZSGeExNCHp3iHjsGv/JMK8cG1SVOv22MMiFgjIABjd9bIPbrh0vCUnpW
NfTzHNAM4V6tHvHT5/swnEtsogUKwkma6mCO9H/Nbd5tIKvvqpDL9eHOwWgVo5PSp/d6knWGcoX3
nVCm2OBOXTkIe2Eoz7E/x4wj3j9IRl8MuMKdL6q5ClsD5YqrkGnlL+X8iO0836v84m+vsPlieiml
hUa/Z9x3EY3eGGQVEmkyhKQnN1E3Fr80XBdrdKecj+z2XThC/sxChjKRBEHvf1weuKDEYr8IPxA8
DVMw80K+LAVOMMdzt+90Ke5oKvWnIpitbdktDSCzJakUWYhVa2F2lbiV5+YqHtcueOS/fCXtTo81
B4SVF1PZvjOX3gD9Y0a6Ivm/maVccG/Fe8tduXPfbeyV316zIysU8pxvCLMKjSJyVmwv7sOKV9oX
dTauagzcR7yXtZikP7OPSaXQ5dSb3D3xU0r4HgIOJTRu1heeEAqjkK77PqQo4lhH5WD5uQWN2Z19
V2gnI8I267Ef915VOn68l8UWBHbe+CiTjiL45rR//OZxi55lmVCQYFpLn6pGjHW5DcttudJAzfQ6
V0W80IR7h335GvGSiltcpBY2YUr+UulN32w30mfiVT2Yt2SrMkx3J6Z0fWdiLo4laUJWCGMF4f/N
MEKdX6lLxLSdA07dRjoBw+xANuTrmZH0NfFh+9pVPAXLqLmBNdub0GZsRIy22tHcjC/aZJmzD5vT
fRPBxPvZsOVUBROjOki1VS+bkdHUmRsX64p8OfzEKx/UDo/GHEWD8QIfm2OS5c3M9Qs7E9yhMb1T
zSWukM5tkMREiRllK+D3kXn6hbHWQNin2baP+TyVNAIXnha2QnPDkfWZC3MhvmpyMrNz2scoFMDm
MsaO3E46y2zuR0xZFK0SZLU9wDFIA8T2hY1yUo+uOcWZbRJuoeviO3KU44CWwgvzWw5n2UR0IRjI
3gerBmSFxnlBLq+YM5l/r6oAwG6Sdvr79ZhBgdcyLuQ+pAurkI2ZXQAVc/wNtvtB+mJYiS+93F1+
PfEMr2fLB+EiyqYHRfJ/qVSVy4VZJY9qY+eIJ0MnAwSBK6Dlo2RPLrB6zCHo1XeWsVs8cnmb0ifi
RnWzPHUyNZEwsXnobdVVZxeZ0rv0xj3Rh2QRVWdNPkNWn53xZZL8wC4Hh3rO92BVySdl+iI6PWi6
7NhK+Toe3CIwkrGpD3BG+FYgtIXCbEZBB12GN3JlE1mLsFzHBnKtszM5wsP2YSV/8/ARIK2MPMHv
E6crabW1tehg4WNkva5oi7/C3z9kHVgfA+Xd1T/CGWz7e05I1+yv2xYFxkfxYA6Mx3+E4jaNNcIw
YgUODThEXZ/6GPuDmbpkZ4PJrDMwbtWq3XoBzj7I4BR1OGBsxUBVbtmC4Dd6UCtlHjAOqi/PQG0G
qHRsRP7WdwwOuKGaMJxNsG89DK2AS7BAXgG+CsgSooHnmpm45yc7RqUcBGYoWl3duPttjnZbit0R
WdrMAA1nNttL+VKWNDSeorvgVn4HE7OixgFPq5BNY4SEEB+hfE8bPPkg512RIkxQ/g/xwJiJ5Sd8
gDvBZgNAZpBKK3RwjzB+mlId4WOdkhc1O4V7Y5bypJwedQSB16Vx38mLjxiBaEC42QuP5o0e3CVN
lHX42t/oYb9/UhcAUqIv6X70bDuvFXupwyJV3Y94fd4VxOMYIA/2J9x3UqrQ1ZHA+kD3PuYIHPuJ
HRBT7fayA/ma7b+hP+aBCHbaNV2RdIpgndfY3TbIPf+XUhcQks7LSXNo3cplLJmnfZYV8pBD1dO2
BpoELpmSnOPAcpI4bytYroVLLcX9MiiWOEYUmB1ReQ5eiiyqaWoRAwwIBuj+2SY2M+6//QMqPuXn
NQiv7To5AEFIooVSLAZlh6paAE6qneMgiHQIlHdCf1VOMdfHHFFl2yFUW1SEdwshdJOZvxbft2Tf
G2tOJ4oS348cnfWBY1dazAAUslp901NElvx7PUHFFcrvVEWR0UlCtPv/8LQ8UKZwMxQ1dd9MeTSo
Eu2nJaB+SXfvCuHjkEVhv/0oqhszawHb4DhJepTZR11Tq+lJLS08iklXTyhMRPgQH+5FXX6OHpo7
5dk+yxqRf1OYKGAgSDwINp+u+T/osCOEsn6b0qrVmUix+udVZej3PsWy4zmE9Tb8LlKVSB+6UoFv
PNgHV1joPf0kudfCb/y26IwWciH2gxU+PFDoh63lDKh77kR+4ORkQeMOgib6AWGyKvrEfNARjBop
zRCd+zr7IHAHOIhWMHAqUaP1oZadtnZSkuo56Oi/YYCp5r6rtRUA4f/BqfEklullJr7J0rdO7UeH
50pQojrn6gvhLP9NI6gnx2psqdIImO1zAPrAtP4XFSXcIvN17EDfmHURe/hIp7ZT/nf2A9Mxj8NG
F4qxXLiOW0LLCPSK4XkcDgIAhEE1roldYvQVMIo1CeXZG1AL5uFOkhG6/MzXkMTIuYxvQBg3jNx2
2k9xd3sn2QUPzChD4KrjyuPQdlUauwR7d47x81poIolBbNzcuyenU4DDFUMunroooJsPKV+/NB2/
gzNZvGCtY4mRcD/cWIRt2fVqrlOjDCHI5ojmUWP4huB9fDKmW/LqMs/7fgRTlwcgUdOKerZmSWaN
Thitlbmo27RxAvj4nt/14lkzrcrOR9ko9Sgew0xHfr/AL//eRurSz9k1M+2N/V+LnGlEu5ygH2P/
VrimgnXBzTI+ralDuMPesvgJLzYFJ8M6t8TH3BXNP9FSb5nUnTYSWrom66XvqkenlR9l0zTYWqUu
lVn+OyBfIcCpnm3+rBqbg3HLzqDSA+P2GQz5kl9p0Q1UEw7lFwiQd4zst2Jq7KghK5LDSYV4TBds
lRnvQNRhUPKWa+po7iFLGMlgOusBD/lHc8AU5BsnmXC2sh084a9T5bnNCFfVyD7HevGQrKpm9xfW
9x7UIomnlfgMyDeWbWPTZzDgWdyYOFHAtVHASMzYMOSX+FJ4JwwUZ1k8rrknaffuZZQIB5bgNSO4
mKke8JH2dWedLvyDW7PurcRlCQSfmg6Z0t2Lo0gmiyibKEmMtvmW0eEi3pQvgSXYJPyjx4xd2tJY
PExRHJkIeKe4srhsJw07oixcyGp1yzx5TurrR8o/NIzqyJ0VlZ8u9stOugXMDWEz6Rxiza6lDIay
e+qzpmEzoU3WHD00i+YlMyFq122rFUaV0+eTqF/B4Rb4fTsMwprRcT/4lRI7KSBFO9diNT9tV8Zg
u+464jyg8nVx+r1mXnFFThgAncKYZCHic/mhTmZDXfBzIgTk/KQfjHbNpQ54eTGwDVkVj1Osk56T
ISeF1kQYIsHUCskgBV8HeNyoRwI14ACLurVXNuWRCnXbv24r3NEvb04dXKRZNCi5+NgaE74PCRrU
ZbzZaBkffIev4Vq7hWnUknto2v9W9aGFozBSPKXDm6uevf9OGxIMxsAjYxowHxHecIP6m5mpPcre
NnsoymxdhWY5BMaYzsiN7cBwjAQ3gN9cWDj826UuDd4oHea4Xrw7UvdWInjCWx9+GdD3GstKG9A5
vQPk3CmZrc4oK67N3g+FStOR6HAQYC9wa+E3dVfTQr0ZPJNO4yDkB1VC2G9Kkbbfe6e4xs6cPEsL
45pda1nIvvai2gqk5P4i/SNI8tQIs6h+g9u8WYqseMCGiC1oypmsnLwlyZrwhgJVT+FgRGARGX8u
YWsb4O+mb+aE9ii+zyRoPVest8y4mZU9UZnD2wKO0WvVhCAmG2c53bpCW1y2RDO0ZMg/CoQ2C2Tx
6OXVObzlpxzdIjVuQiHSpYOuBHv/LijT5U6z8b02t/KJ3bQO4882wLqaHlpm2eQhkFzNm1nKEtr5
7J3rMueSuYarFabb7JnexWSguaqmCbsRaLODMdCOJWLva4+NT40Vp+53KkvYHNxkhQFCpARCulOm
poe1sQbBf6SwvGz60gWeVFOByoD6EOaTQLmeYb2NAieGXn9H6A+HKafCwtd72cwR0HWft7Ky0Jl4
9sNbFLeN/KtIaLGBKWqhaGtbaaxfpa7qc6nZE9QZ0CpgOnYFYn9IfcnVHHv7qIimPTOv9dfHtZno
9+WeTLHXAU47dxMHND3soJFNRto6w3YWp+R92UUTkjR+HhEZKCPc6S1RY8D7XXpqHri0iPsBp2CE
FDGRNDRec1PQxeZqZiDp89Hfe3b4TRhabjcWw2UO3SZhM8bmLzSskO38PFVSLEV3X4fbkjX6uxp8
R0JvVHlPPYwzOJgv/0bpgaA/0TFnbNtwMk+AV8TGBQE+kYA8wcdE078+NsnYILCBBiKaXBCCcd1v
a/88j8RWqsV5GB3UxI925JgHkl53wQvpPLAc3gXlFOi2DHQtRW5RRtRZl0OZGylbTfg7g/ka1jUx
8NvxC8oKuF1ZCWWOHwncqhAVWJd9IWlArZboqKekTiM7jAzovCKwBN7D6TpPit6YwGVKGUloVC+5
1TY+BESRjmri1fgxVLXv9v/QEuhVUIdwaYYx2wTQVcMLZTXgtnO37WpNnvrkTF9jzM1aNCxd+s+X
BWlxh4g5v1tR2gcgNeFm3EXfHx7pCzXf5qHY2lkk9zysTCF4j2wjteF2d165Y29tGZIsaCGOT04Q
iDFdgjh7iYRtDCJ23WIq/I4TfI0SYLGnf6gQsr8S7w83dr/fyuiy7SJEeDb+ZZSEvGvQwNq/VJ+F
1HfgQb/7DdSRNTL0mv8axo/euPqKf1H3UO/YHYrjhLjL9qGo6HuwXvV6D8G5hOyXnw7O6X0HcDQl
xesEPj06TG+i9Lw35zsp3xLROJdRhqhhsTsYudL8St+dgppix0Ex96c991dX/M8wMZFwZXM84s4f
35fmbrdSo9ogR4dEEcTGij9UaXD8nV3lFmkkHdapO5HVsBecGOH51ZXn+pLxU9N6dKbsCIp5hsi4
ononJ6Ds/mQXkBd8eYLBUJfHYUqGhgvsWLSYi+IrIzTWMJfb6EibL/XewivkSHu4UVA0ojfQ8UBx
p/7p8cs5W2LchZN0FceHPHpj+qA9YHFh6a7h49Nazn+cPSOZQhVCsvhN0Ml7EavCEcN4jEOFSFWz
KgDKn3juJnv7UUkz3YUwTamSjV2GWgAmDe4Xc8lLTsoi9YU6o3XwQjZl4sAkn1SHlm5F+wYjunQw
H0ZX7tbAktxwfwSpWajcR1mOPZYilrHKDuIakpSt97D7a4LPNkZhdO4pNy3vDt2VE6u7DD3r1JQz
yVvfwEaE4WVdtrKu0QikzyD/5dBllvpg1VXFcwx5zoxuD4FUaXWFsJP8v4ceHNEwcjg19OSvWxaK
QYTgGgHSajvFMsMnYFJV4ObUT44nDUfZuZ93kAVQXeYxm7YvGA1qh4ycawNo+2lKRTZo87EH/hWU
f3j+m/NPI9MoL3V2Vcd0SY2NuRmMDHGMhnB21JPn0qwrJHkI0EOY7qkt4S8/S/mYNzlgCTLOk9F2
qIbEP24/IRN10E+uuGVP2jDWWO7oxl82Qs+Fftpogzg0PkCCZMPqyl2kEcrw9+rkHxcgCASQXsgr
EceQBnUcObN+YbnPZdLx82Mc3D/7mipakuMc5VCK9kwqgO15sL5DcVzl/z30Bh/RXW5I3wwlpt04
OmOpcDOs92uxgG1+8qXOoHaPdR9CjDXUz2of6V5O2t6kCHJgDfyB5/5kNFgKTkavtl3mfg8yUue8
lerkkKYJ+16QosrgbAFwVih2i9bw6W8cw7y9Yl0umJgG3jviq+ShnXJrYnxB3mDiNpTTyziu4JWJ
TamLvBdssFAOlKDrkOgnmLA4bT3w0Y2eRqWm4Qna/kZzDAosxJFrhZEvp+5S79jAC7hbM3ADZ3h7
Jkm5JAdJiQiCPmO4DeHi8lN3kuxPcC7EP5HmV5x85txO+ezh1Mz7KUmSOMKVshWl3Yjq9vYFHguB
DfgMVaCplYqZ90twhgPoS2gL5DrioEs5bgW5hTxi8TXSgR2okriIrRZ5l2yeAlK+bWbi+d/81x0d
owiOlda3ha+a2PMpSZ2sXFzwvb1pplm6cDOVuFVgTj0sSAE+f4YSWUh/M179ugWqEiVAkTlilooU
FrkI3qsnWVFC+H72m6WRB+cTSSo7BJiG5CDkjX4XRf0Gtw8i0zsLPhJDfxHcCogKsLkZpscePo7/
69Kx6oV6mvdMrqoUnFR/YtQxr6rzLKrsDG5/8XrCsRqZTg5AUym67YO3kkNq5FJYY0/ObM3Midtu
+LMa5yIPWkOyanqw5MNCaMYo9XANz8sHba8fozJOhYDFJDGoqgrn1/ZLJA4AznafKurabeVHMn3b
IWf+P4Iv78G+nzpWd4zsdr5YrGafgG33CMSJ1EadM+v9yd50035kDBah2blGaCXzgiAgBz9aNK9a
g5cjkigoMFXeZDu6FlqyRZrWYDx4lG9Sys3BEUirw+dAOvCoVwjj6KnwQHDdmgCVljDVV3x5+LFv
wHsJr/fN0BISn2G0uv/07lWwlxNlmSiQrfjzJYj8OeAkHrYPQQbIvtxrsZP8PomvpUVMKfQGFLxB
foZCrCTJ+pdou/twZE6s6jYYW59pYcRfgjU57HECqPAMfuDWutxUrNmeBb1v5batWSqhztN64Tf+
ydGV5giLj04Ynw1OSiRUju0cuc9z3wxbjk99U0YF7Hj4KUq/3G0TN4s3hRYYv+uwq5X107rbFTHr
Xglf+anQfPxFF6zBdmXFPKHbTDX/cwMu+XeLravXKQ3ofrK25Hvh7VF+jhrwovJtn+JYV14A4lH9
EADhwKUgJMwoMUmTifATsNYNsnJwCNj7dNp8NGyehuHxkKpNUGG06yb+u3uxKdg1eDMaXB1rYLNv
AYEdF5cyWjCHzEr95arl+zE6Feb9QHdt/t+e1Ht3mMAj8yYWgbEeUjqsQIVOFRUxtHBkP7INH8Xa
3wbm8Q0SN6V9nUn2YD1hTadbNWLIO8y81ZjV4PYIp0UzAqjPL5cURn3LOXoqbkxvoAq+/l+mavWv
ELUKLx2NosH+3ZQ42dSpEdp2L8v1Wlncs4NP5Aw9Qs0e6b5kIxktvYl+FhqxPqr6b1ep2QQ6gahW
gJ9/+EZfSxgVq3HvI2G/YUdGp7VvEo1k4pQIiROuZXOmsLLSc3wAkfObR7Ey5VfiQ0xEJY3eXOkZ
ClYhTxb/hLAqd6sqEfGbtnbBOyVJMmaTGn99nXBsmf+QTRuZvqo1SRUgXSkxjiu6/cjJKdVG/J8A
qGZGhIuWwLHzmxZxEN38lIxd/lE/995KL72AAg7RZLgePNag4UX8SLe2wDuK2oMVDNBzX9lcmzz6
mnYXJHFTJtNfF1vXl1lKuELaWgzwXSHvWrFm4k/EG8KlZMmDqJepKPZ8GuujV71iGZiFaj5DRiPv
l+nlhQYzgtUQLHMkAspDeH3+6GbysEyL+4am50FNW1ifvr4itPDakrQMkR7wYWSfIWCad/AgAeZc
Wa4l2CXAulmXWsnQtRa8ZKBdNUtmBeQpL3f2HrVl3l+12TI9QlwSz41tT/mvayvULJtONrduLpbo
D5XXGd/K7m9GCqs9RtQuOdC5GcJf4f+7tgeZT5zISMNz3QRPS59PclSHWxdLCYhNKv9vWRxa/leU
3O1zFJyRp2CudIiZWCTdjaT4yGelBVmVmljzSI0jbXWsboDf1g3shBlPN27Fr6EYjjwIgQURSrzS
9hqkfJuohup6CrHiLvDdQ4t6xzh7mClUIYa/vQT7Ys3sEKwn0glShYa7xp7H/tounBG5a0Iu+qGx
F9FEjZEWA9TKBwD94KV4CVuWYCyXeprF8xhoEc6yyX5Gj4I898tlHZwLjSlipm/nshar/vnboWDw
GTKB5xC40kEcryNFCArTjPJ0oDQ9cwem8AYcHxFOtdgQotyxtFfGqvzV3w5oz/8oaC+HSLMS62Xj
DuTqPLvyoC186cDEWjAjD0woWpG3yigXX1BWNtbCMAAEUh0Owma7m1FdsrW+IAxI3Yo/aQNgBo6u
y57njHYJ5SFrOsRNeQrjl0i2fBtHAOjygNkmwbl9eUcAe+baWvj6hb4jc+fSJxM8OhTMveeqSHmg
OYOWj9zHL1kpAaKpBfMCP+B7sAwySzCkTWCKqEIjpTdKMY2ZAe03E3ZPwYXUn5/OgVTWxjlJFdTa
NOqxZeOSBUiYsywy9LH+t8HnMsQf3YvT6jt02C+N72Ehp4dukcw0ayg31CO36f1NZvEqmrZUE8HN
Uh5VsBtxc4YQN7TBo4eXJ0e+zRimrjGX5xw+nA8O4G3aecVLQF3gKdDQLcf+l3Kp9nAS8Vy4AGo3
CpVCHfgu2MPOqOeIzgqfX5C2TAtCKEnsMFGckIBq2T9XRgz3w4+k/IVCmWtFqFVjKVa/5YqJT5MF
SOYhIEJcPgrX/Xqy9GP9imAqMDZdeX/CTkElWkRgKXyNKw+cfkJK2bZSixhl9jui+28IhfoM98Se
BkDuPMKlpimoyYHfDX5yhyN+jGID1XF1/LbISpbZOb9cc6IGr3+k3tPc4B1VEwMe3t53Y0KsxLyU
MFhZ9CrWUUhjkTrTJTUt14eqccH59nNXGLpcjBcOKRGy++UbhUt5AK8zCt/ez4O/y1bTC/kMXi7i
PO4C4A0o62oAbfDvnNTCLrUcfYiBcRlPM+4RY3btTRqLJ0iVEtcmgEKmPgIyFro9IM0MxK6TlAFS
7gl5fuWpqMlfv94lgCBFwkSK15ztvbfzF10VgYF5M6j2HBdy/HdUGP/bPiqI+kbBmzj4srD5V6Up
OsfMHJdjedpzXqO199tpt97TjlEgvs4+t0aJkFgUNTiWJxo4ucFWBxItfXrbMuVpKQJXkSSA2ics
IPexWlbvkU+E/R9Up6JcmFJ+lYvTY1hM/u43FKzB75WqEHfqs1x+XuX2EMWnlSxgbrAKRM3UbvQI
nfXvx+TcPiuolus1f+6VB4MsPjpGH8zWF7Dek/MPx69fJK/SgOgppM+Obb0CfMArU8bcx6A7WBLA
j5V57txgBzP0fxt5D5RSIQd28wi26LotSMxiZcyZ5gud5cMrpy2MDHM8fsGCtmZcpshwCCaQJlKb
wh+8hNRk98Pkk7btcacZ2V4If1GJULe4r9i69P9IFI6NBMLu7+jNLzlnXeau3veHphS5Pcpyflj3
zXWVFqQy6Mq9oNVcOD3cuUDjN7ufL4lW/u0D76upuYaoREAdH0WR8/NFr3VNx0mAafdSmKyO0T1d
9Gv6Md35qf/1oulCI5VQnuykZQVSFRYQCd2i1tSJXa7fnHcn5eYodDHSu0NFstNOCzbh9dyKCqDj
l/kvGulXTXRNe7G6tLv0tz7lcAHuwNSWkKbm7io70rUuoK/5jQxUbd9ufoiaIPgwqeGydI70RNwA
cEiHkWTWtXxjHoUfAyI35J55Rx9BQ8xchm7QbqErkzyixiebLA2/db9iRAC46xqPQcdqxbB5IsZi
iVv3S7nQVcpdK8LBB5pYXvZvBv4nU+ZUUQpP+mAmz6uj0yhxsHfH28lqsRHcGq/jHmSAMpoX7Klr
vrB9BVWO0sk15g6QXwx7tEnqD0uCcI0sz/CRvwtzd+C0K8qcpynWZ+qYbIchzyAtOpop9ze8CZTc
CmQ6OLV6skmWHym0fy8JbkSmix+7d7LvgQg/G/bVwC89XbOHknrA3bQiKSckQpyknqhSy+/nVn0T
thUcsODPjJxKi7DJ/J9RRYa6p6DP2+eBcn+90/6SLHaxy64cx65nQa4ji7TXr/KnYo0OYVxODTZf
HUpGN6dekc1gWRisD4k/697jd8g1S6ziO/6lwV0nqiU+uLREatbusvXzrwyb5z2NiL6Ck/29xnLa
L0aIVNQMVbhPSh+u9dCVLGbNsQlyaZyVlVhPcdKviY31bRV10RbtuCm5QiM9GMGDB1xDCfPJpTto
DrmKCSmGPZwkrj3enRy4c6sXKwmc5zwTRAjE6EuCJYISn5WdKDRiCbZoQvJYeY8R75nO4OTNa6q9
JTt/fa4lDyb8gvkRK7ne3UNLBGMsCo0g6zRrPxGnHdELArZ40FFX8Ig5Kf5dN3pnwNdd1QFNoisb
OapDL9JYLRwb68E6KWYshSOEP/M4oJYqSTocnGSx/0dewZ3Muk1xBvQQadM+EjpVym5sPNLnK3Nj
umOfwOBITsUIDPyHF1F3kCTPLrAZaUD57bOINVYgQHvz/i3f7O8f37sBJkJD+JhPfw66THnQj0zd
9S40ihDsmRKKjEF9rBfdFXRoqyiV3vGCKEJaZUrMnCeN9QZb76TH9lkB3S9NdGqfD0MJR/UjPGGc
o04S9Jddzhdh5d6A/AXRItXJquiPN+7mWDEGA1+Lb3F0JerMKykQdYmtgrt/0AxJRxpbDUJxnu0k
LGMaoUHoF2lWG+EPe1v/j0zcruGt3PenH+3Dlaa+xGDVdjRO47b/hpvun5QZ01OhAhW65tf8aEmn
RD//jRQ09UjmTyFxBL/7+R8VWZ112VjioKgiSn07BSM9e3vvINaSJQvZX0zpKXQ9jiK+tmIpR0RF
bvaOxD4lWFUhVVAJ/0luwn+DFFfi6Lki/qOkbJ3ptlK3F+2NQ5ovebdeBL+XYv+b3TekorVcFCKx
UFdoXqhkXTgIm6Pggu9AUp3mWa1MxpM/YymtpmSz95BXQZ45CVD0Hyg6d6IedvEJVeowooT0FuMT
vfC/fJf+i8/JG7HC12Kckou9Z+hefwyHXduPlpHVtRk5W9splHEq6XWLNFGmfResvAZFUUSf65bt
I3KcgUrD76RW3zyMQ+0K9UzyAuN/qgSSvu5GXQCRI+LKKnQZvRZcdC6Rjc+vDVuAfvRXiWwWfzIJ
3+3RuP5691IHL82rQpsqjL6CbRUXAKwBC3AUU1AxzB1psxEGmf6uUkwpWyWBtzc4M+jag5yeoK0T
YbpF9PNrXCGhAsF28UQwj9A2XRVQ6yEJdINvex54A0vEPpu9jI04M7H1C2KVg3emvAPyozhk/3VT
sVQrq90H2+OFzBaKK/FCpzdRl0BgIfQ/OqiFFixphJOy6S4fKDFyDa74UeUOBESK6vJTEKcSw+MC
VVW+x86lRj3zV5HC9xGgdCk0aHQw6mDjxsMRgygfSov8Z6ngB/Hofp2tXq6zUj8E2joEOgw48r9F
VnukUvh2dA7VFAx+oVykTLnXzh1EpEHSVzo1OIKMvOrqY3Ld1lwtbq9XnShM75Q8NPb9w3fFhPqJ
JcWu0QAyBikoQnfLBKJUCQy3dDt1Oj6j+KqSVefAgURi4v6JccTbPtgbv7W7QvWIpwsXeBNW93Y0
USN8CAI2cvAuCiYVnwzg6s/jw7B+On2nx59BA9LLp1KTPGLBw/8s5Qwcunh659vB3YXqNRSyd1D/
WWmeufzUoT3W0KYNlfn+udZyATNMbEUDjlZWtRHhaa7ekQVLGZFIwRBt0AtRaeMv2MArosPsMZBj
Vk4HikWuQnpjEL/avpCN7Jb14uamENus30+ajNUbe8zT6317BTMV9xcXZHKXCeD/ZvtVFtQU1Srg
oM7g7vnEaEXYSa02VDBTlFv6IsuBitpXI5755/iE2vboKPXNyGJ5XJ4+VQrzk6DXaAqTYyquGYRl
GB8RVLLCpdwg3ZxDtaSgN1dx2tFxRa+UURzNzL1e2pG9WZQNYimMoCOJNWNXACTr3YcLtAjLa/K/
bL1s+YETaVZPcLc0lJ45QsL3PXloTDG+t0kM9mDcEI/UdfcxHuapNAdJ8CpRLViai9N2EM9Mrh28
Qv5bdsEciGSWwF/kDGN2ytK3qKtF9sy3f7J5NjQ4Bk8OUyEgu/7tNgb3oYlhvYc9PRT0FBE0cFxt
lD/7u7aZbc+aSlFDLaoZnBaNx7ItMb+bA9hFXsye2wy9mbYtv5U8IhLBOMThUkea1N6X/eBcbmhY
jwTth3n+KEkeg2vUm6/MJPIWLV0s/gcPFhxZY9b4OF/0z8JVUQ6jOLhqA57tYp3phU3qenbJmiOY
675bzJyvcqUjcrGQRsWI2ej0UbdKIASOxVXgUNVd4xsRBTy5ovV64xilvPCyC5txZUaBus2bHVMM
3NeiQoUgWaJY+kPRO48WXeJftZsiE3/xQmgVwffzQFczVsylxQmUfEs54gIQ+V0RTqHGSOoj2TpU
KBHbjiycWTl1ILHicQ1co4Wta+4NvpV+P6HreCA58p36UeBbSHSIiF+OOa0xYOcZXEt7Lu8aZMNI
U+IrvsWgyGtpm11oo+0fMlJUMVNIrjEyARrgKZ1CxYr0DWeKAPvse/b8zzRngproEO6p8CRUf5J4
GEBl+vHiTpo/h5Mz3x/gIKWfLbpRTcn5zcnIhTuKP+/jA3cV9yzw0mEmEOtYoewaXVM2/xcL27Id
AkQQnSMebUN4uXmdTMTWgAeSOej3X1pfJNu/7sTHJWw7ZjrK27SnxvmivZFw0yHo15VuMMyh/WFO
mNAyBx39ZXBKbmVxmsw2hWYFWVtrmOzIau+IGgzN+jDXmXkqfObdg4atY9wh75LT60hKpsC/v/o2
+jbdJy9PFXipNJqUocCA3rsJYbczwP1g+nqk8GdbzrCPdL4z2UpG2HYGaYGKa8+kaw+yfzg+cNio
j4aWRklZy250+lQPw/UedbqgFTKcRhtwtKZRO1aKlL3h6sN4Oi3wJmNDlw25Hpi+1gP+7aLZ/AXl
KKUcqT4dBn40/MoF4BQvnjQCesvwZ5aIyCI/ymCZr2Lz2QaUHmTfgKS0I4jBTZw4Pb/UwttW8qM/
FhveqVXh+yISdIGJvm6ky0yoFbS5Il81dAtMFMm90QNu78CXACXn2rFu4sJJuSPhxSHbakM5jurI
1gVJCCweCDihQBcrAUaCbbbnFI+eYmsIxlQjlm78vhQTghC+NdF83XkVFwaoNvu1csskedM9Ys46
apZUMiDKBP1Qnpbu+aWAU6AMob+hYsekTkpD0idnmlbcfT9PJ7FnltpBrkRrPz6ewwx48to5QZCG
dt1q+PsaqHb6dFuq+qPvCFEKJGLkdppeZR2RIZyS1B7Q3/D2x9kKJ20fE6L/yvrmg7of/bdtzAY2
vt+iVAyiT1XrvfW0kw1yoo69+DuJUiFa0zqWFlXtxFGfh5uBU6Wcx6BRq8D87u4QgF/5NV3SIRyn
yy1XgLUpdlG+8hjhtqZAbFyQoK2f/NgmDf7n/qKZAqd0S5vS+/Q1kgK0VZWL0AgWdAdSze4+fzKZ
qDyvnY0qCSfJTtjGEvyhjJIJbbiiGqC3Op56ps6sjf7MW1h6ATTxfECnX9XAT9FfEUAS5iMGlXIv
cqlmIOySO1PYv44o2ltDM4NGgKLBeuTGUtuu9ULn8Xs89oROV8/y+diMAPz5bkaoeem+qZPwR5cn
dRfBNXueJhHsxilcDLcNYaxABuZ/D9ibcBYMbH+8eKmYvWh3j81Gdv+fF1ZXPTVJcvJMwjbTcbti
rvzBuftpZOurp8tDhTuc1m+KiZfOCmYL3piOOTXe2V7aznysqv29JRYz6RiPGHii/Zn1Av+rggdo
WUJHJpyQGvYdhFRAu+3GTigaIQsbH/NYXi2P/5In3VN8D4+Ty7d58EM3om8gcIFCVg0AEK8fF44k
rpxNq2NKDdtnMOYggLuhl3NJ3s1D9TVV4dsPe87vD5AmhXQ/Pui1nQVRkFxAM6+vB1lgEWM0GjM5
UCmyARtZR9kRFWu+flCb+cbpbyrUt3gBf/1AtAprc7TD7jP/RAZR8E6XFBWTLZy58Indx5pvNnvw
+pDyVQmxrEaH1OoRFHpO4I4QN9RMHYbQJN6yMn/ak7Y/2nOH6cbrr8nCV4tRPQq4yWjDJLovT3Sw
CfOTM3JwzK4yxtIaj83c+aFxvtIu3VgNo1+jcrVPvyW1MIjOPUrSqFfx1kwgttsYI7EZYPQ0jKww
iu4zn6eqFVmx3+9VZpleb7bS2kXyfema42k9JrfdffGbs/Ig3eW1ysKmWJFNdPFsndzb23JyGGVg
m+SA2GlmGTpiMbcRlNhJXXbCOOIJZ0wD4otRxI2r1Zt4YLuuT9OVY/CXV/r3YNOVoYXen/LHFWEU
drIaVvb7fEk+O48VllAWlASpQOPvbC0J0U+Df0ZPpUZJn7wS3Vl2bSmh6pR37iy1YogPNLnSdSM/
a77UhJzCgV4f5s3UBHkKNa8m+WyN2tA1EudJX5Wa3mpnUf5cTYLM9+RgyfgCLcn+B6xV2ct/oGeY
hl7SIY6Udp4mBlCka3Pb9SxhlFUZKBYglPWBLntw43dOBFZKBjaCCWKijOk5EJlqTb8+BnQV+r3I
Y4E5xiYTwZulQy/E3ms6BVB1tJJNslN+qB1t9Y+jgXz05tLkQsRznpp0mbZm80iW8lx4n9TpGKAE
//mRxdBeNQ1ffuhJqPNHJEHOLmeFVIYff8O8O0tsC6mjMld9dOnfkXLpvHty1tD46+lDhZl3fzL6
GfNGv5a/IbTmtSDQaFjUxIMeRIjH/dfmtO3JO1wQmCLkOVNz04pNouDuaR1ZpYha8BVufsj6gaiV
LayptA0yrFKtKqnr2wxM1dQR6hh4+A4QpxVg11BqO4JTmExsT1z/j57ABs62g+PObFv9vmIwqgxy
W1psaeyMVWV6sWTBdIr22kn4jdGjioe3bLUM7SibvCaNmyTBRP2yxnaPKUmBQ1rCUVPFM/w+vcta
TClhLF/i2t3rVf9VYAT7q0fv7k7hOlwKoOwVVZOVu9UF1u1Fj5LQjPkbiJrXgFXriHVGB64X5ma1
2tznQNhO8UAdKhJf8tQttWP6J4rRtCLHrFHH7j+AzxK4Kb9M2p/4mdTbWPjCdVgtbh8PrXUfQ13H
LYiRvWRsnpW6PPf5Fdn+YKZVGKTAMJXx5hLdB5GkGSoisx4CqPDgjrqk1KH3I9B64XOWTlSLFRcE
ladSI5Yj6WEpbSN1q8DjSl4cgVfN3un2U9vBxx3QYkym2VYAM5MexAKbvOGsD/GFYGkxOFLjdygd
Sj6ZQl8dkE3RNHNy+EVVZME4dUTaRTcIeyEAFY3PbGMXkdZCS+3/J46e2JWrBtsxqfQQs43prOcU
tv1aMPtohUNh5vR7y36tTr2BHHinAfeMivRmgXgXrIoWkViKUKi4dVi+34UmvV577yBL+M7jwFO3
r5tkpx/7fbBcxHZ3AbR5H2OMtY5WMAZtO4X3x5t6910QzfGIaB+7hDEYxHrDZWd73KHqMSYrDpRE
QbW/nvcPvJGGMvztIwJlT/WRDVqRqKCbpzX8ru/pc1v6XBVwoa0NV9VxWylnlZwz4HA9OjBphDd+
cwdaktZ1qD3qjjGHJX8VW08VAqbQFp1lnaggANm1nDUENYM42c4gM+0y1z0TJ3I3VpQjoc00uvyq
E5aOkfJD6MHqcVEelqpacIu+jQY+gmVKuzX9KDs3q4wS1hgsNOo9nUcpgbOVfGrK9cRc7X7y12Ne
cKMNtN5LNugr5Dhiz7UmrnvLAPevm1y5DlRnygenSDMXzHQCc4kGSdd2vJbVxyF0n7dCJfUvRhZK
xupQB2y5J5mvyud/tV8C5ti0SvFPWLE3v9j6tdadZ7iZyTuVFZtaz70PhWMjvQKuzAl0P9BGAmPc
wsj0F+yU+cxo1B3fSVyoB2jFIbxX5tgMWSkiAmhZpzVF3RzhJ/K5Px2LCXqf+4mtZZ0y6myr+Wag
bgM9PQj0Vob1qsoJna77Dig9W6ibyLWNOUeHYwEGjkPikDQqU0YFTeWeUssoXZ3CxaLTQXtpdSJ1
LnwXZ+nXs9y4+MFn79Wru85r46rZt/ldUpgAhS1dp8crBJ0/WqXekA4EwVhX9DFVLcIEj7SLrucD
MxFeaIzTeeuTs+jncI7+Hv5OxEXezlASI2Zx5o0mmQflrzJJ3eoCyblzGeZYxhHO2lZaPHBcu7GI
t20G6IeyhXpICUnLojObouXCwyZiigJVSxTR5Y393kQTDC7NhtXqEe9wq+cAMMqyYN/YQYrO57YF
bq2b7b+Q7opuFiYaelDuN8IkC0WXmu8RStQZhBPIZ1Xs14CMtiuQkdKubH4oCqlmYxMy1R41XDcO
JSIB01SFY1FL0JSP1uzyJDhpg7WeTi6qmnIQjwEolQ8l5104V1Ka/86A7wHycDhJ44En7FO1+u2p
yKa26E422qRQbK23RauLx3dJ/bbHZqRoAk8SgnqaIH5AQ95W/J+B7SOsLTTBnmNh4IAlzdrbJ5p4
VSr07eqfEei+vbYGii7YjZvT0mUV/jKLyNwCeNiZ0Zf7r4a6NhbV7tO3XAKzWFGh+BSY/qPnVTZ1
lTbtckpBBfCkB1M97BJbQpZbepezxx+z1nYb2a+VhjnPce3d29Lz6nsDzdlkC8nOAFiH7AoGT8zK
LMSzl9Dhj2/F80Nd5HUsF5Wieb6gJoD+NFxgAXCs3g08ZpT0tvwMFFN4Fj/Bnn5kZzjgX74g2wIH
2BFaT/xACYyx2YNahQRLizOSVtC7rSnS/QzkW3yKFbTCm/OcO4ndo30VR+FSHqtTtleQ/O0vqPL8
eYjDJkIZTQDe3OgenBZL0IZx+VJpBhSNisb7pBASm/rwMGdOdlPq1m4mFFVXZ4JPj4WRQ8K1mXY1
DH3Zh7CUw0bqsqpis/GvDpR8Lxj2Xo9l86aJ34c32f5s6va4nq+9NDKH7iKOp7GyAIxPr4uFCtOr
qVid7K4dBfF2uFU/xD524Duw65CSh0i7JRDxLsU75O5VUV/wuBVz27vxL489LcG3SGpaSVK4PKnI
pAytXn6hKz6mpz/90wns7EBByuY8IqFCDcSnjnyRr1RC37tRtLPUN3zyZZYsbF+dLIWSCsl3jBY9
FPCkYbCKO1qlKZqnLy+ByTqpBUw6WMe1/xsIv8diMLV/GFN0JIx/4NPaRg+OaoOqTdKEiN6XDNxt
IqkYQUp6daL+I4teJAX+PTiYoqmkH+34epFTEikmExq5soAM6wUjG7zYeiUS6srlPbNOfi/+abnN
Q3CVf+r6Pc+zkOhqZI0P/vkO8hTytt5sdJPN3fNI/18p/nt7tfFGLVaPIh+CtbhWtoCvMMXEEOb5
iZ66FcvrGAPzY4kjVw+GMjoyJ738IGz+JYuw1oVJAJ14+9wHtVVOzofA2X7L7maRgm73svE3uCPo
KpXrOXP4vnGpm9am9pbG10oQvR3au/iCcKk98kGjDs7NTm26PuTvcqaKVwRpW9lBIkrrjGFCqaw6
7cOXYfxXFOxasaXjRLM+46stkiSGkNqLObIyl3d7w432NlYRLCZ3TE/uxVzHRkDxlzMUuskDSvSU
D6GIh6tFQ1wRA3k4FHinlYhT1P7N/zu168zP/NVbM00sm9mZh+aPoswSe92+mVxz0BL2h2f8KDvj
WdgVecurZhNfvnhgdDwrGD6GlSKNQUCnC7XbljJLwLanxg88fTy58U/c89vm8Dllm9Np6hfVjOuN
4qOhtDGpCacSAhqVuPsgdYVK90LkyKNN0e/iDGpf8iKyyUKiKBBJGUPjT4esvUP8RsyABWnp2SUt
1WCgkdcvTITB9aT9YU8r5N4cHW4KKRpBKyokBuG0YeKX9vUbG7khyBXprBYCi3Zs8cMkg+ZXXLxC
ib0WY5v9NISRIjX5V9rmxMTTOz1ZmsIF07B0SJhj1FIl2cQn3+jjDWhsgmdTKUp13nSinl9CKP5J
+WVyUAAzMcaJB+UGzYj2CSXuKR6/PP1epjnte1NkZTnD3LuQJEUMMulgW/COllJCxQEdW+Y0ETv7
DpWSrzsM25msxzlBmdDE4IqypGnd6wAPsgxwccrSmvnZLf/q7ELxbelCala7NJQP5EEB+GeRNpqA
bx5ubIHsVJnFL5cwPx3LKs3BwLhYvhg4kwxpluNdU1Gw7nGcoiDWhrx0VRFvKdfaD6PZgA4XaUO0
5/v8lUcPAxubZ4BQXAKQK+cOOZ0PQrn6V/pCvkzlI9aXa3Kb5IRUUs4zAW7gBR+ivok8jmSaVSIO
AuSeXHhLdyuDsaqc4EilKkRsZvLnrVgV/NhTu+Ee2WF4gjKljDnS0iCLOPf8YQZ7E4lic/ngD5gX
MhUvRDKMHf5GR9ktvqlVJE+wWXRAdFfRX9KugFSHZbNV04JC0qlEuA9V3+2EWDUUd17KynemDcas
8H/nxD7gbG2Hi4FSBvKY+hpBFq0XizCQeQmKxnYpJkuvKmWRCkRXqIth5ipyMqW03k9r//4YIUru
BI4im2cgXYzwXn0CKRNl80yA3uZ8AcNtzo9/7hwNydBbZ1BYqISGJrVVqTa4koQmyfLGXPwhYjoS
UeXbfg0kbkHARGdaemzPDZwV6Zs1OLr5raYZ46VtH4Qm+GP6jE+qBiyLv4Hh4ZHJU//bG6QjKqnS
FaJclqf5zWmvoZdObmHfw616q1VghJIX2BAeWu35Js10/lCL6zjKN6V5u7N++m7aU9xhdfintSHb
3woes5GLycSAhR2NKDAeEaaNN0cH0n1tKxKi6gNFHymNhUgEu5rYWjR5czB49XTDKuYXi7IArEGx
Go/ShGlJB2WxicphWX+KhX/VB9y7hHOt3DbUZ9WmzigZez/VBR9PG/LwTNOfmnXoyxR9vES1g5o5
um+WzuSo6wpyHcKxiJSpwNWqnlzQClmSwB6mmhP7lbQLG/jA1p89GZVK2e8iKJQ3TnHUwD4HlICG
9Az8lXjKYZXkVJauII8b319IJXN2jxPhB3stNPL6ozeX9wP2hW7+me84UeQ0J48e2S4ET77EkuST
uoxSV/NItydEHQXcnR5VbMb8/wKMu1DI8oZGGkE9sDZ/IPct51oohOIotvbr5vSWYonkTk5DBasN
nTBRO63dxbHHs56eDHhnHEbSY5epoXE6SUfbsVnEdMuTr7mnIp+nZuVIkd6lp8/tpwqHonZ9siJh
3KKTImwJpCvAl9hF1sf3ox4XvUfz7h7l12RKTfuxH767oUnv76Y9/LcIXao0rl4DSbGD2/LI0qmm
A0rnf2jzGuWAhao5MsAKiHsSMpIqcAOUYB9SbAkJzxsByALOGBoQYx11X1VrSGCh/zzPEMKBk5HG
KfFHoYyFuPgmeKwOWRIv0Iu+WFrkVg4l0cp6e4wZ/bVn67xGANfeJL2hx3VfSulBe6Ys3bw8n3tf
9jeBOOQPXzmWQquJavPa5C014Flw5EKNpbqbhC6paExh5L8SiBAO8O28BbXegHB6B2cN/k2mb9vF
WLoxIXiaR/zAz0Xka9ohV5Z3SPCReGZGAYd7wD+nnb6INBFV+fMLW8bs8vhHoVOnOgAzNTGJ6HTw
l+HGLP+t08z5uhl9oJ1yla+MU7xU9Ik9LmqU7EqXgdqJGtxfuRnE1KoqaoltA8QGg/SVW0ctx+2M
gi4+KSquMhBMZSsGaG+qnPemMYaIwvVQnsiu+nGTKRlH32KVEgiez8a0rRDtNWrMLLPwQVdxAL93
UqSSw5xnzxhC0Q8bnbi9Lh8kkrqhr7n7Wk6hSaqYbsdbbDQX+sU0sNm3buSHiE7koXld9abNG6y0
7veP0XJhAzqIG4/Syyk76LRNmjmuc8YX0YKs0BA4B51zR565RwMiPTAWfC11hEKKyKBCGIPCv2aV
Mcc44j5u8IvdOsTOOG8XjK1rHv7fe23/bXYTxrj+PhK2CsOCswNxZrlWL6mZV/8CQSDkWoRspaHr
eHBBN7UeUR1LDeqhsr8Gc2EL0rZfDVz3G03o210+L/wtaFuxZuGnhLSw43mRY+IMsGwg5rKhrmra
IKEkYsMtp8SXLcyCfYgsgjp1XmR4m5+1P+8twlF4ppBPjXGrn4PuVn1rPwRK41ggkplO+2z2lTfV
yMyA1ojDln9NrzNocM4IYKbDZZfY5/tFOlLNnmNinXz0KhK11QrVEaTOCGAPRkEtqBQd3IBTGekD
GWYhgc1Ijc7ohkZiodzD/2EtN7l171YqZ0o/XQv0iZTk0sXvxs5bfSbEfvdNeNPm0QFDoNj+nKTS
mOTMkw/OJUaG0+K6Btih/2TBZFl9IxEy2AlNNIEzzK9+XNh1rttL8csLmVKTrfFv7ZVymSZu3bS7
Ap6UGMGf0USnlpDPahAC4rkJDY8cYlPr2F6C889xRdjr/kCQ8nvmLLZmmA++YvCItJpP95+GB2qJ
VuxWpEvVqeXPYm2lQdkyBkBCR6n5nY3yF8XEDzqBxtQEcTjynXt3pEFvSKiAgaJiolPyCS7H9oUa
iWRMpA/bu3WnxVmB0bXANyG7Gitib2n8ADOeVGAExSwnhzz/B0N9nRnfLR3mRS4zrYxEJFRUXiyf
Ohhhjc/JWqfks1yhjwwt0/g0TUSV6gjxk0XlLegkZSCq+gUipZBfX7aMJr7CYUPP6S0Jge7/0Y61
2xdQWF+AwFNdSGgx2csUTFzVEtXtvnzc3+eGyZvT+7jY4BTUyBNZxiVOjpoyS/AfYhth+OpbhWvc
DRO1uevqJvuXVb2tB2NEwJGsWo7U/Z7o/S5YZGky0nqcfGAiGPNNdKctZucOu7GI9q/fZeJ3RGiH
hUs0jmyyz54lkuG4SRgsYgtKH6KirlEgbj8mowXsbfYudtp9X4xVIidCOPms05DxofxftvmUnitN
aKnT7YgbyEw8P+7yFqKAishLLpsss+PYixSdk7gx/S9f48osG3VZBpclmld5q9XYOi7uQtYyq3M3
OibJawZIYANNKsIdfexzoywjxdYJTfgfBQz40Yd04QKCj6fHtal6gkVKvdDVMFa9hrZyOaxPsmGR
5zE51dTKqSv4qyt443M1QMa6t+oiq8NM2k6V9nGhQF/UYZyzfon8b8D89eU0N4Y1BZ8noGRd0SCi
4tRECDZHzdgfiEVQ0HXOkiWROpOgIoHeRl+cK7GkaySZ063de5mamkK4/fgpYT20AAlYD4yLGxPm
5TkIiLQgOzK4f90K6zs+jskVAVuGuJkmBNIXJikH3DyOa2lJJHl22n6a0AH8vOwYlWO93ImOcoe6
Hboemkl9EweQqbLKuV6dMUXmzS3kcBNNGjrQl2gZXodMfDKJifRqObI05m6hk9tiD6t6r8Zyp5X1
HdkzgrpITfOvTu+Nx5eYxIZa5c8bHInLuy0Mcchu7jAnw5De2hxuSzQaoNfT/oZi0k2IQol9qQ69
eYk+581Rn1m315aE+9YuCmjk97KVOuT0PgdUHLGvfVESiuFiqXGolEmdvtK226wyY/8YNp95xUSK
YKV/mhuoO/o9jO8YoJbEUqeTkl5QTzDRcE/fYoThUTScaYnRxkUK56sVMKxZfmKs7H+3y+wiHJhd
wqcRl8MIDfg3XVnhegl3H1XP+fKIdF4J9GuaCSr18UpKx8td33Mae7o5T5HAuqq0IeJI6SyV7N3x
xOmwAWWt6gK2gWvL0roCDbiKwjkE8PRkfdLY/vGZRiRwbTQ2gxr1hYc8xZxkJzT9/NFu4Gts5MDK
bKjK6tiK6OTfzzNPXfT73swA8lXHSiGeU7b3WDKbiXfzsadAVmKIfxcNiUOP19rC5YAjFkqEKEgK
mMBYp33+d5DKhSpgvh7NfRYs++26PAVABJ+iJdh+fooSNm8KxsgYGsRhdZ70huOc3BgCgSCKdZpo
C11knRgeQ7Ug0yE2GStMVO7FNe/8ijU1ZXEeR+uwIpB4pw8zY6L1Toh8O/8s+cvsU1/Q4U7q7L/m
ygwXqosZ5VTDpBgA+rkIHSQ5BG/oQfYZXcsVcc4bj0ZgLBdkgTx5UMKo24Jl10+rJhVVsHhMzVLK
CdLXbeHychIxU7nGuAj9uGshSbzYnS4G7XWRWsDVDVe7c7sUTnIvuJLCdImRJszaP/aD5LyDEMfs
taWgA2qVbbE5+fis2LAV3yc8RYJWzo5AwPYIiZIHNSBJoJ0lPxA4Kyx/AUKg7jjLqho759eQ1bWf
GEh7iQ/8NieOE2nUe00bmBV1/OyWNBlhWMWFIDXl7G1PVsR5+4b/Ri0XkBqXsx7EnqeLY+OAywb/
43v75MDoV2/fgCprtaBMv6dD6aUseVTQR5Ifot12ebwy7VK2ImCgUzMhr3+jOcom5wgn6gRzvHOX
ktJuH+IX9fNp1LTazEMBC28rmjt+T0BBlVDVmAb+fFOuTTfT0gHf7XGugTngUbSqtPjraz2cG3yF
3jTRahdXLQZ+2HOXD/H4CaA+7Kpwy+oyZrAXP5+p3iSle/QrQC2dn/rQlbGA2Hbtx9xhYbK9frVJ
UVqmOFo0goteYhNGL+oWZDBNKG0SSwHlGSLpAt4z1DKCSAtxGm8ZPwP1GUO6/7lZXOgIgHOyBVS9
ofHCdE/kdguxFzs1YPWDDHmPo4b2e2AphDoGXFmmL5fyAGgVA0ouRG5w+vq/F8UgBpSznM78GT8l
+J84UhNaPrQYr8cWXkfofe5q1QH/fUAdAI0N8Jg1VQQW74S06iJ3X9DpHLpmYXjo3gRN4huy+mYd
UbB1FbyVpHPtGLX6r7kJMWLL/4tu2ZE4MUEoeG8H7/OjFeU7MXHuQq1GUsWM5FPtCTpY7fAlHTrR
feLPC3L01EUMpofwSx6KYrzSg9/9QlqPdKLllKSEb/hwY3tk4F/2RQl2gSKV4DKzxyC94LsuEJcK
XKoHqt4iNlpZUqXXEhV0K2ozqUd+WluvGxNURObOQKNghEIafWA/vpqTQ4k4rhKgJ5ihQe5aG4+7
H+x6lTjkyym+wLgiRQclGp6fgimqARwUT8/3paQPlXhWZHX5dua5yF9aZeP22blFr+93PmjAQwq8
YPEhjnWbodtAioXVtR+DimN0fCEXqY53xh0I5K+9OWebBP7+ZJ0zmwknvPNjBQW3U50BSa6HaoeW
Lulig6bxinj2hHRy3drbZZ8lAIs7FPLaoxxQIpb6bDl4GDoZZrQX0abLSDhbTqyS2ww+andM3MhD
vyG9Ru3FhUEBtKvmA3Ac2DutmywVyfVvRW9KYC+OQr/VDAYzsH9IUeM0bLxMLHPOOdeUPAeBMscF
eQ45rQNKXVbelUFGFRt/j4lQBP6BEZ/JJGHRwsbDX+x0mmC+KQeZ6hTDUjlu8y4K8AGk8QSXrYj8
5uMLt3LGsSknYP2Rb0Cfxqa4t/OxP+Eu92XdFT73ZjbcuBQhuD+lSu98e5yjD3GG5gAlbN7AR/lD
xqLgjhM/12vFXu7uBajt4huZEBZijlaQfVJ6Grw0Z5KKWUW2aCWNT3IN/iUdp5F+UJR2KV4i0/zS
xDW9ejcrbm/7c8aD60KD/Illi+5Rzri5HTU8pvkyi+bEPlc3p+lWXiebTv9fovGen1dxlg6eWcVF
jMy353qAA6yO47nq/Cl9VlWsfp26EDAJMxggRhIYiWDtd8Bygao0QoJf3fCHWrQeZQ5m7FEZSld4
0ztW3OEUzSTXejhpgXy3/i14G86NCgsc9xsHrVRVL6xMM3RKrRPv08C4O3U0G1cP4Ks/25Y/MLle
dW0lg0l3TOId0U+IdWk9qKPOy9t5qBYgBQX29+mzJOHUYTpwT+wm/vlsEYORueGWMTDgaAAq3+oF
FrqxhosWwwHdx12VJR80EvawaR/XBUSuwkcMR/O/29ymU8mhDqlSb8EWrGe2bknDK6q58ez3vxDF
mPU1Inhqyaku6ni/k2QCoXBheL4RAUn7xJhp1ZcxhtBg1CTZ5+M5ElmjDqWezzXh6Z0f6qbElnhn
W5mOcj1YLvwn7ZDPPYW/f47iUR9QptQVigikUWBP7mxJWvv0Rc+D51Q1bzdUb8gVil5sp3GqRhiG
AQVZbsm0TsOtpHLON/XEKYZsTTDEWsfu72dcTNcBO1O+DyJoijnLFc4MCFs54KopGbFDgJEn49ux
hSOpDYqk0mxInowuNCOyIlo814KUBQyBG4dDGJGuq2diIsALDoTGGSCd2jxvor81cHB34CbYv1+1
KJSfgR8z7/xsPSU5aT3z5iMMRYO1Bq30oiXh/PFM5GczN83O3gHAnIL38NFjxcaVn4S6ase/ck16
JmpJUFaga0ZykxK82JZGTdM42xcdnmiKkYQvo26C4yMDivpiJshvaoLVqn8lRb2hedlKX4otG7UV
Ei3Q34JSko+sCmt9zKicnmFC9ghckXcM+Z09QV3netpMAMZPypnG2nSpenZOafLKTueBZ8xdjj2M
BzI8bKqDsFiZgjw0MuMRgwOQ8gikUlMNz+T8Mqu+sHx4XGv+aVez4icqWMYVrt7btYVVg6QIHOg5
QONVY8ZL7eveLYZNqyRvN5QGmIjd7mW8TOgcjLj80a9H48k2rlFj7NtIjGUWBwL4s1E5QHrHmD1E
0LzO6AIHwSsVY8qLQVcPF2r061VC99ks7ODPVtRD2YXQKdIzbyMTpObV/WbzGLhrmLbDbYBB+aoO
JVTdNuqYDDANF97Lk4Z5gfwbJRr5/Ow70+1F1xqa5fQ4Q/Jo1R0S9574wx51Ig4cnphMZ7+NI3T6
7ldVwDmSONTzhDBP5dOB28Wg7f9ACy73wuyIWki7uDjgpZIHhizu3z4jPgObEoy1vL5/LRxVNWcI
TVF7P9zjOzJTZ3DSKhyJQ7c12EbwhrJxiuLZx5L9U53Pepuu0xF+PJhSUOLjvRjjGPNsNWIeAATA
L/v6EoaUcbkPTlKqODnBn5PXjnoAxqqOChQiuJTTBNttVlJrsbtYeWFjhq8Up7VAXpY0XFGx+uva
JNzaEgevuQufEqvq4uKr6IOilW+qjt8oXjI6IfYHec41RbYh/CqjrsPmnqp+aTXO/askVYjcBJUO
KbiO3bVdYMIUqho8zKc/PLffr8iYWvReW6np/uhvKcCiHWqTYgA3PZxbknjqTXy7TuOIRWHIiLAJ
mEC0xSvKtriKDNcmBCMnYKI8UiCV1RcQeP2uplwu/4aMurOEvzb2ijZxvfEgLPfE/RR1tE2tAAb3
nvTv4mrI3+kfF2kmqk4GS3bDd2GyIr8HrF9LTPwhuFDRZuQVCZEl1LuqwCZpTws2P5CGNwpvyqPX
VH9UI9s1GqUfDJUNLTN7iDmCnslaHH9CQHJg0if1jjx6+1CFavgqxe76Ry+nXBi5+KeKKPbxGWma
8V6Ih3Ch23fQwB435wINI0cETgKwfB5sOe0eZ04QMTT7LvuclnoNzQ9NKIt9YbMQJqQZC9L48P99
3BMCBCaVIKXw/usmJkbp2Nhu/0/fuhzD3PwApPKStbXcaSr3LwuKXxTG79qOYfklIwUsBIkAj5M7
mNRLeXZXLEo2F8iCBugD92n8DYrGTrFBkt8C1AbCb6FoNVOVy1NLWHmAE5QVjC32mxXT+I37+m2T
4qMfC2gu+NxOWYiXK3ZNuEEJbzQXfR9s2hTMFuiRlKIP3ZJ+xDR0GEb7k3JTwvlyFMF3321i/OhT
qTDn4qeyhdQ2CN7dBg1x/1l/HbEy4jzDt38ugLzAtULxJQrGpHyr+EfWEYSq0mF2xpO3g+Lj1DiN
ToefaykwHp626gupMvmSi3zUQRxhv5q3+ZUIR4pBj3Yyic0YIRAIXIJ/WMDU/g/5fn7spfzOKEjv
Knp81syj8D9+KjV98d3f0YTaLhHLWAmP0YqU7gCARz+9psFcjEcOO/5EpGI7kHQUY0KoRBfrNNnq
sIHHiQuNfuklaKdq/ia8acWMP8UsyPYws00pclrn7ADjm0vTr/L1ZkgKxukoZDoWE1jG8U2O+8LT
/2q5nityCGN0BaH9KtVusujyg0MZPg79UH59zC/VyXlJxLXbicq1USbxK8WP5/lDNfJPOwAqxa/B
0Gfgr98Gb3vR30njY2Rb5R6pAyPfA3lLDgbzJJgYL+9zDpU7D70OfmWkAK7x64zDhv5QKa0N2bQd
/LyssYBrNgMumci+uAwwUSHDKkw8QtXxI5rSZwceyAC9gz/6BOoaI1STV2Lo6ysV7zWr4HFLqm7Q
gINPR4Gghx3KpRkffDahxf+gEDEgwDiQSkiV4UxfR/28i1fffOvA/uMGG2xxECaRvBGlzeAr/uXh
RNrru1Z23RpOKqIrciz5aQKD2Q9hWw2urSjX4Yopj2Q5vzUMado+C2uT4dSQVT6LvP786TKLUsmA
Fl9KqujrtEQhGnj1BWDf0qTEMd4EUHOKGpvluEZypHYocKs7/sIsEyWQwXvdZNpN7s4pMELBOabc
mNDcwzxv5mleRlVN7kYbIAOFoTVtZ9JQpXE4ac0xEJ0EtM6W6C3LqThc6yoV4p6/wCT48zAvv3bh
EFu47p0jd7llSR9AICexMa1qykcLIpjlBoS9GL6I4xExPgaKatCMaolfQg5UVu8HVuXDvjIn8pAg
V7UkjIhDpowpqvOhYa5c3y6uaZN0dMgqQepeVFpu6YMjz6IOg4bPPFd6QKCc/05ZWl3W8fC4/BSL
3oLCzadcg+hUCaH/jDDSgrh5Yehm4zyoyUwoo8NsJWULgm2/puxS9w1vafRUZ4k53YuRogtwKSOS
99X/i/woazD/h4dSt0VnVtfcz2gakEjsV+Xp24AycW4m0qQnjjkT2rlRYXZ9uXhtkavq8NlL6/RJ
7u9fzBFEnuJHJ8nZrjJFDqG/pnY9lAvF/Fn3/rw1K+X2qvcN91j2yYwy/YZ40CefA7tOcHfR1ZX+
baqTq11yhlu/2GkxY01mcRqvE0bPXARgVKo5IDPew1W/nilDt5bKH5bikVxWxDoPzHL2fS4K8IaE
ryZCwEPpXNNurbJFLQt4RDUQSNzCU+YsoFDUYYgXJz/7qKgRV1mXka5QP3x8mOWHOZamJgLrr8yU
ZaAJDyT9AwRSU84vtkhySIrjjQxyiuRlwiyuwnj08lW0AXKA99IopVrdPvTn5JupEcHsLlF1YMbi
QufAwGThPwToiq61Ga/gu26nBshQteXZ5pplxWZw9RSmizfFYK34A1hRIgthXMqodvM1s5/VAaSw
n0wKApM/X2Ye/5mToi8GEEWzJ9isAnx0OecBeAsun2NteT70OBE8xJNSTdZKLPeTYu0cb1MezAKk
x9AHYuIeulp3pZVrGAw/WdI5ASFPEVxQt3N6fWt4nPBs5vB/tgiktyJ2vljaKSyzD8HG9sqHIaOH
itQ116nhbXGG2u4lhVj7HyLCvHkcit7okmskiUWiADgLUXPAbCK7iEdg50kezCY+iMaCUxLPKHQK
6GhdZzzFurGsCvHK+SZn91HCbI17D0pylF51w8d0pmhbdxAUQmseeq7TXZfxJhGqhffh2p0JEQNu
pS7klM9UjjAGK/khNpzlAScWryFVN+AvtegAhxQ8oNDYZwov+8d7eTtzuiSWbrkdOjGbrR8o7z45
eUMYxUBjj45/OD4WyFYNVjgmJ8iDMdrwOXKQWvc04stVzVLCEDht8xOtvLMuW7iMjQPOpJuwCqX+
1SdQRqxo53DuRcrltEk2G2ZwRUyhoAiDpAiBIbDuauy/5BAkdwOYwhMwwuzLiQm9aFogRAZDxMLE
U61DWQOtOM/cl3pBvMmHLxFXBv80jDiHGkaEHz1q7V5Sw901qedOF+vZ64t920yyyi7vsvmRRwNb
ej1nbgux4BhC59UWJ6bXm4vhq+N+VzxbyDcxPTnixe7pLRnfmYQhQl7pdY+lVN9hdA9GtjZuoY7O
RNEqfZXYaAWY7hYNEGhJ9bLW0XSlLZ+LmRxjwuesNDUm9mh8dQj9TVjeIT8iZK4cc+F2mD2mHWh1
6xvFfVXEabxMLphxFU06c6zXss07zJLAIRzo7l0PlBs3RugBICkLIDD3ROpOTgvQTVb4gCbRk8uN
5kcVFbk8d1HbVoEr27uzXXazTzgJ7s6bWYOQ8wK7cN2MlkkuizdUiOVnhx+uBzNpUN7wBFWpf7AZ
FwEfmWvEoDFeWwYScUM+YHTvHvmEEeqeDcZZt+dyvi2cwnIEPGaBXciduhBgS/XBzi9b2hYtd0Bc
hvSjhIJiV72gCR60WkSJ1kRjDwVgQy6DCYsxouqP44BMhwNu/gyMUpsJqNg96MER5S0H3KvfpqWX
om9aAjiSe7KHG0Fm2khwHdIurQiO2Pfm7C5iSxZMoOWMoAtQhvcHwIl0MIP9usIiJxpVCnif7buy
K6myEXMkqiNJ/8I1Ojo/frUR04j7Cyr5GyUt+/SSGHCg7HwUn80LC2MDVrAvHRBz82sI4txwa0SR
LC8L0/YaXmWGA6SPM2IJ3jsUIBHyNA0CTO6b3z4UrfpQjUTAH2JP2BeellCf1wFnbr8qA+zOz1b+
02Jt+FS4LGHNDgTRO+cEQsUli4HrxztvKnJkCdKJtae1RpggKhFTS1fYl7WnZ4XZz0/UCE+llJea
nM8ZtUrO2dJnGU28yHQ93kJ1/e3PtXUIUQMwdsyYylYob3c6RkAkjJ+b83yK8pMvda/Grukv3Ywk
snIo9THqF6vQBAJPNfvadP91bhDoXIySJ/6LP4Mhrk2zBwA527iNNkQ1cbX+63nDHSoF5esAJ+1g
HKpETGJpGvuI8VMRedTMBE3AYSnrqUXF2RvpCX7ppvb4btcxhFqm/BEoytR6mMpMAI9+pjYps8eZ
C61tjlL5xQSK06SG4XIG5reylY2JwnrrqJ/Lolb3Zawq0A7f/cZZ/9TpG1Wc3EXPpa/xS+KsXHNx
CNmp8EudqEE5oniNJJT6BCUVPyNGtADZ9FKIHzctmW2PQG/7jPSTn0VW4+q7dcjihkeK2dU52gl4
NJpXg04hJQBw7vGozQGThR8GhwmS++zkGpi0jLVmg7YU8r5zkADmhgUM3nlMlXoqEt4HW5r+HIRB
MUm6xvm+qke0GxhVvx8+h9aTzlIiQKjzY8WTufB+xvUTGeFvb6gNmRs3OZiA2DiI3okrcw7uesTh
lya2uJdrKKihrhjwtHU/MU/Iyanu6Y1fnCPt9jRLRAC30IUeSYOBr71msmX7orVHdcTJI2nLRl3k
1wLcK/EVLpFuAuLU8DI/GA8N50uAm8+8a3IW3qvmQkFGPyttehjPD1M+20HmI6RpSXU0k1pLQoSr
fyxkixYMiktLkgRC+u2CTiLTT8nTgm7nc2Rj1kv0GfWrFdnzwoemyjsn7s2yrFTpPLeZyjAksm3f
CV46pUc43yCMk9anSSFk8juh9qrJJWJ8WYWMOaWUxlKJ76kvqtM5NUadFNvG9kvm8G6oEx4xg5kI
gWQ1yiqInpvzXRdG4ksbb5lUtKXXGADUyQl7fw7DoZYvEKOnszfFuxecZ+eGBNeOjwEc7nYExd/5
b6w7vfr8N8GbjErBJgjL/zlaa2JLb4olGg3yLRMcZn6V3Clm8qTyHD2WC48yc113aOGNEzwkxlrG
03kMS+1TAYic53jBc3iYQ/E8y8Fkf+FD2BckpaWr4Ecrt5luBdoYVrW7pI745sHGohyu71/k0LgO
kUxyDwEFTb+aYm58KIHODnRuFn/vdmwUqltm3fdx3ARCxtAmt8Anxkj+Q+x46x4TAbOLeCowzTLv
OppUMuVUyzcgEJncn2YHY/EmnJwM/Q8RR8mhGw8bWZXz1r6X6h11hRMghtartGu8fRmwbKVpIAP/
tO4yggynuIXHIhyqut3CkEMUMoe2i2jNRicIabXgk81YrYOcbSWmfq3KssamjdSkQrB1UeccvtJ2
+2EQZXQ6hzxkXmCYlzi8yvGcRe/9WOyN4ebV3WH/V9vSV398DLEEg5lpCc1u8mheEEzO7Q33+lXJ
jJs5+KjZIKw+5Vq2caySEX4/1ccppnzw9Yhhy2zWYkOlxafTTsH408WQ3Kpa3lTBiZBylr7/bfZ9
0+i4UAUqZdyvpzJkG/TY/InSedelIXmJJpoKbB9xWeOkH0XGjspuvSaKqJ7XiB+hlECUeelJeJb+
YPbY0uoy2HV8OapPnBJaRCHBADnFwgmOMv6FksVqmaWsYhTU02b/zSVVcJEo8cSjK6k/ER8f88zF
vebez7NgmUqtdopS+x/9zH/yEBPPo9Sfdf4n3Zy1ACwjYOkbdlUS/FS9iZuL3NP1EjggTFipIXQN
9vGfiJyay/fZ1gTb7jq+TGU2wNjXcNISF6TxL5BbKIDDVA+Uq0ZozkhPFHuriHnsv6xVJ7Ad0F3H
/ys9mCUMd9QRcWuYlPHh4uOD4Cgk4HFfPR29m10D4TePzgv3LopMl3DhgOOkSroYXpcb/qvgq4Bl
CfRn11HN71pzFIPTv60EgQJMTcrdeob97znFfhqQIgSbQeeLUt2FPGzMcc4U3vQ14VQP9B/+uhzE
tYtFZPL4YOJya1z+XLBjVAs32C2hT8DPbsYb112TiyKhQY/ZduT1ou/iE4G6f4C/w3UzAsqcU6eU
lDSfA0BHJHVWYNwKz0aT+wvNCVz2oFtVMgNKu4zP/Y2JAYrFZi2bf7h5p9b/SeWuh2BN1dGJRRGq
xrvfBsmanK1vtBbXJ0d9sPTjPoF891RhmXV1Wbr6GkSmYtA5oVPz/HH1N4bEus52owC/GtYFEfeW
LKnfbUrg/PAC7yJRRCKx+QnHuQQVpcE3vboVwLM7ev04vLGROrcoE7hrStfOkPrpPMsBJ/CXIg0w
YAZCkjZfpHRTzPjQJHXcHPQuqeVx6X9RC2q18ttCdH3Mh4oCGwrQie7YFXvHMYk9CYdv6w+kqzhT
mecK1bUair7BzhVXn64KWHMlcZrgKt/8clPPQ/BIF13L/HsMZVZhno6ZVtE9i8QSXHwbK9dk1Ym+
rMJUJFEaT1CVhtTfpMW7fRFYU8hSAsEUVG+OrcND67TQymniIGCX2mhpb9ucElVm0S0lZAzz+zyI
/sFdmBGnOP3okPcioDjc/hCZNP4y1njmEayzlhowk2HIUydhQn+yT/tqxa+WkQTiIBd9zYwC4X6j
d1i+dRug0xQsIepotxX8bjzd0G1XJ7vKYVgQi1H4pr08OitNtj2HI+mTcn/jOgwgqz9E7nPNSfSq
o1gI09ZM5kPRDyn0DZtw0aOFnIQjHShiq9MOcuIxdqBJUkXziVlJp4fERgqI8wZ6Lr4Bt5vtBdpk
VJYo2gaHevUkyVCzyVH3046z2J6aVGeuktjw8vxaxAPZkNv/QemCMvceBq8xGjxSjy/yg85lWywz
4NHwraAblkmAEqDbtaUgmK0vUrGsSLm6C+y4nu8yropukps3nfMZG0qSAuNP5CIlZGqPrevgZ7zZ
0W8E3AOrcjDu5TOjb8EJCTs6b2VJHu6uB/Zz5SnhPHLCRqdaJyx3nu1RovEFleu79/MGvZ9RtzPI
r3vLmWadSc550hi83jDC2Socsa3toJqaLmye7YslPrFAoHNoyzQu/IEaFskf4LsoBToW21DqkSfa
wIgpYcJaWOYuL4HZ32iJsGRG1QHgX7FpisYeL3+SgNy0BwE2tgXCS5sEByoAeW3Cr8PnzJJZqPom
2fs6QxAKU4xTbJEYGcD5ISjRLUBEcm3J+4VQOX/5VIGb0lQU6CK1PkhqyJCEl3ZOM2vOD65NrEGc
RX04euX6TgU8qGYRBesEpEv9Yxme9lAG0aMsG/qdajCgwe04BwvmFSuatcOcRzWOEwIJjDXgKfY1
2MvvV/+ifdpxZOY2c5JMFJs5F7+BMTAsv4z04hKXsLY09bcakyl7vZO6UjGsUWwB4Fx0b0ZOuIOn
JRVtWBV7XLteZok5ujycaqRAFyyZ+6HJzHrTBvNDjbrUr+aANvsSiUjnqJfKOLtaQz7N2DKr6Gtv
FVXXpFl/znOFVOIezsr9jBVVxUMA+Flh1FE7ILZE2e+KNSoxmCG1HdCbNOFtrJkFsDBLUhk4dlqD
8TWhs5FOlSKWavysTd91YRJidmjtbu5VQrSvMb3PrNlEhwdxQhYXOBeuqIzuWPjbfF2KPXpXmfYm
tktHIrAxFXdChKr8tm4fUeZ5gR/1AK75YkO4uasl2N9aXZ8sRf2YDkHaNBvid7fX5ii3Bpotz0yj
00ip+fKIkDiw9/z8iFKCxZqr5zQ7blk80AVBRKI5vism0zqiYfDA5fcgpkgZRd43wSNVva9lNN6u
IipJKCmC2b9S5Pa/BnHRR834ettn5BsDH4tGifEBPRnEEbBGgSGv/1Wdenp0mU5Wz7yX8R9qt7SG
qLrtVtdOlWTlp9JcgLO31KiHnXvOgzr1oe+DYwRKG7h9qGJ9oCVb3q6/ZZZjeOIiUvKQGzZoF0hP
pjWB0tlZlswDX/AjFhITFnRKKTwrpRANRy6au4nNjqkK2E7JRN8L5zm6KvoxnVngUJC1FgQhBa4y
EFyMjcL98dl6JizravXXFxNZsocak//QBe31SDRNj0uBXjdSxMgOWPxZZHmJrnWPWGM7hXPrkk1A
hLryRP3zKl/NEfZ48lBSuAZtsj8QYEnIvl/C09JnWsOqvp+BXD67Qf/3Fmlffq5amrjRrIX0kvx1
HvDBKzeEEufg1qv9UlKbTbAb/ZYvK2HsoYAN+Zt5kOFZkoStd/rs1cX1RSXe4V1p2ZO53BqDD0ms
kd/Yc/qJEo3gxePGyQTmqf/SrLWpqyEzyuP047zIzovu5B4+XGn23z8BkCQVLQuJJiraFpKtRdTm
9MQdjkSDHPzlE0uc4LNQDHrIyyowbMa9JdxIwLhe73ztQDsMbudXfUDaqtiSCkIC/eWinzT50MNm
X7x7fjEv9rH2Orukd427d7pm8czHKUFZhev9fcUlkQPLOH1sK32nwL3sz1HS1z3xZVysQXHgH/86
fKWU+ZqLzeb2KkpCC2wZgw09Fc+BRfglATDJ34v3GnjcSuQFSfttY4sp2DomrzyZ+U3B2KxxgmDZ
4MsDffszpwX2SY6Ep3DA8mVjKpbSHZ4NRuFeazIGI/lvAbCYEgelZKMAel6IQjiAtjwrH46uAMZt
0CyFG6UWZhihKy3CCIuN6RDWlJ9vu+qr+Ho503U9GTmTi+SlL56MDAso+9GL9hRMGf9ZVWrQffRL
24bzevJOwp7RlyKHCBHmkQVfPT2EeUMNupKkuLmgM8Bh7mwokP05k1H2t6f8CqWZCY17YiOKjFgJ
UweD5DOFlOOKdN8SLyFovr6GSOLuOr99bmRvV/i9NgOID4fZskHh05YdYz8chZHKSaWtjM3xo3iO
rlcJb5GYXpmpFbRpCE66DJtGEgy4wYQPnRwC1WtkvdJ5zCdQq05MrUiKPw/6lrB2SlYP21SpIp/3
sIiptad2OHB8xsJCja5i2KBaY+/R0GS0t7c5FbhEipScMITAdDVBccaBU3Tl1wcGr8qoIlz4Y7Kw
hRfii1Li56tBLgfmZF1GOxtN8GzHdxcMknNQUKhKD0sVW2680Cw2J26lP+t2d0vnaq0QKPmnTt4m
vUS6Hr+zl1ypX+hSW02oA88lKsV7/68BdGl44Hl3+Bkgdhg+1iIl6AvmDeJ06r6Gt5xE4ic4cLQn
82N6rgilCCG4MR/PdnsMABDwsM67UNfqK28c3exRM7xHzCyn3jN8n6yDVgX3mEIwr9Yb5gFow8MB
t5u465CrQmmCVH+MM62Ibeo7Ar9Y4sumzsjnxTYJ8yX7r76h2iOqtDZotVcJRWpRdPktbZLekwuE
vykZmO4KfB6IqOfpruYIp2kadrQRs6YSoBth9thG9JkIRvsmjz+2jIJjHtvFAw0jZZVo963cFter
MKbi/UaX1C4PUatepDxy6NphBpR3TcKWZPcks5Ja15hsxv4V9MFaKQgWW1k2d493qmfrG9J2Bck/
uNzik6yjbUKkyuAeSvpeJQa5l2F8BzC7DwIHsR3hbc3JBTJomlpodAsCelU4Zs7qf1QVlyh0BzyZ
3hx4uliWMS+30GxkkuMK0GyO/7npe/rM0CMbmGdgGVL2vcWjEWy1X0eRIbEN08jaBP5SKEXKMFct
AJK/peJsAmzIPeLSEJ8ny0V2jX1U5QdGTVxMdaTBJokdyGA8NFzZMwpf0mdDazOhJ/Xe5mex6fzF
E/pJCsnR4jaK/DV2KgPb8iyY5a3ge+fC9cwX+WIVtwGVJc7UqkLbYUe3qS0PNZWafLbcPeH1llWK
cxthh4tMU6gXKR0fJmQET0IruSfINqKZ8mjf1TH4nSqcJsEsvcwxi7X6YpBSnr+tKP/yC+eWmRX0
6Csyxi6xqWNzu1WKSnWCTBzWy18w2nH8snP3nW0WYS0OLIGMkP+IGt49mjiMb16IKUWAASeEGgK6
F//LZH0nzjLlFCjP20KwKa71vo6P5d4Ugmk+ZaEF7Z/CYuziZbJlwXSPukSGBFTT678Mgrim9tn6
PKwNguf59TYGvjbFurbhJos24gIP89jnSYZkavhy8lhpoIX+3Nc+fmqC2fm85C2/uD4kdg9S5v3Y
hHDpingNn0wNbAm2x79Y26YJqU3FBTKncK6DE3cIy3HoRYeAb7HYuM9iLmicrHSGfhoul9zl+hdZ
1xZ4NiH4Yir3og2kosBUIMgEJrpN9euT/7qDFOu76l8v7N0QeGhxYrjyoJyW0ZD/m3aJunn1fhqB
GhieIK0xnmXB3t1t8/tLDqJc1FEUUobTinE3tfY1H9SDbjlBAeoLWdVxwsbLDOohPZReSE1iCmm2
pQeSdH8Hj8ndxw+hVJdVwuyPNZb0IqBJ8i3LW5COdJkEEtsUeCtKmh8k0q7T869L5pNUzTWzS8Dv
/F/k3oIQwKOVomEN2SFdSgKFq1L3fx34+/jtNbn8ZscHJjoQLwGbUc4AqJ6bPSZJn+mEaHfIOEjr
7ScQhfO9IBIeO00Mtayd4wk4ml9HFuWQY1/Cv+kd7+k2uoBvurwVMqM+gV90qAUOh8ZMFftd2yQj
kfKK7B3rc0D+mgcwNb2VGh358sP37vx3pO36EiK2gcuyn+HkSwVAf0Jn8kt3iIlUBvqW0iw+JfzP
Yfd4x0GPfECASm52BK7+NvAv9xCpSQY0bCB1kNhQFTRMJjRzMlTZMXTyCgMn2aByJuSsYIBKagCs
Rj8bcUTpK8sy9kEzrkr8HYw7AsQOVERepm9hBJoNi8hGtqn3hYLAt1UIzV83EW8yIEcaXOODdZCV
rUheLgpg2KWle3Ys7SEZCswNpjFB2pEeuJi0MzFGVnLMqL3jZs6AJGt+78N54Th2wI/0PuG47WcL
/BQVkPi25nuw+fym1q7meD+LmwyvV0eKx+qvs0tZsjuyKOES+m1Qps8gZjA1B2gWQj6caKlrFWPB
7xnl8j5c17qNHr1QmcH4VVCZ/fRWsprth/ImlznDrtJmwdtGLTv8Wh9gadF7Xq3pWEyqXs2qes/Y
6KRKmqEWY/GHHCPWs13N6nlz3WUCD6hNrvWU8uzUlTqxMeD/SpWx9Hqv8Tlk9Xmf6QQ1QU3b1rCv
Ie2qeXsQCHIDmgZOgoTvIpNm0lykz5ySoLHDpxYz1jFZP54S6haWUZoaVN7lSbGanpOVIZoKlGkg
IjdNjIJzzpRJkLAOgUzWnZOqVkrDvubG5iVPG2aZUZE+Xjx+EaQdyF1R6YC7hJHjzyLWnyqfCJdc
Kh3CxuG53cLEE3mNe0whzh4V14N2RFNWeVk5ujrw5bU1K6lvGFmD5D7jQqExZWuWDHeRjXbahtWO
Efr9ZWofcK49U8/6Q2ZOWNKY/FqF56uziyc//97Rkz0zkF41nkTk3blPCyMa8g0qNNSpm+qCMxwi
eS2EsACNH22si+I+tkzI/q7hR3MlaRVg5ZIxjTuhOPhAwhvak2nepulgLZUHZ12fg5xKL4c7WnLm
OBsmzYrgTrvZFVhuMUVcUtnfeEpb3uiucuFSmq2UMudibSvw+5pncOQVaJqOqrXhu7a1ltyaqaDD
Q113khzN52IazYG/lWgx+39jSrcUBNABm7n2dHZ4hRTtvYC2wWcjILU7cQEfxyygB8P5c5Buy4Ts
9PW+a8jucfBWCM9u/NVaYzJqVWToVWXOLcS55/E7GLd+Vpct2/WdPD9Rquqc29SQYX7Rg+mPFIs9
fX79CdoH2PcVooTvvE8dVGbXxB7Opw0+v9/0cekeDFRTj/5g1atcn0u4zYxr0tzxNkYh33in1Uki
a6AUoGValMMhlh0ClgEMcIEjZIQcxd/c8l/iV7xrVmzQ5N35xKrFUbaRaUpwUF0vMt5MqjaKLdQM
1F3SBY/mS9JhQkbzbsKXl6i8Q71gTFKGrEc+siWyxkl3doeY2VmEt6GTQL0xbmcyxqNPVeO9xiRJ
NNpm3yTBGlYm1hlV7Gp28t40U7ZKOsbeURjBy0BLW21A5F9suBlZ9BMv8xEY6gf5v8ZyW+m1hLj9
sG7+50F8AQxstuAwrAqIlsNfTYTKzNy9N5dFUdJ36m6tl+3ojyENZTxIdi+jLhR4pscVyF3mp7OK
jXxdKEb6mDk6EgIqy4fcoB7+0Q4tysxTQSLTbWmk7UrrlS8jGDsfEMUj0b8qoL/ZY1xzyPwKmqY4
uBwMDZwTXpX41kF6npP3/xFI2XAht7yzvHL9IjcYKXzmiJSaw6o3vt8nuop4YhMmd9TJ7PguWfSR
pmo4W4PjKK5ZjOHCG36avnlzjEcyJQMwNTUos+aWBB28ht+c+sBIG02wOsMAbAsp8O5rceM0AMO+
kVPWlfxBf/o1xvdcUlj8w9BhKbVed+yYUT1HycHHClp0z1GfoRmFZfZmiUZvlKvHmSH88O3Olz4a
buB6LV00G4it2GyrayVUsv+UaN0b6dSzz9WWPBvyfN7Of0L5B30+HxjhEz/s62rHBphoLiXXpRhM
t88J4EDOgK4zGJe6rHBxbLYFTTF7chkIP41nTGKHsWDtEVwtBrYmIOFYJKkEl5lzhxQmJlb3B1i9
RFDFBwNtvdHY2q1MgNkUWtxyT471mq8O6VH0XmU6d8T0DbM0jrPz7shKC5jrIjvNeEkSov77SmYg
CTPUE3PfCs3p/sDVpPqp6zQq0KikZBKn6WW0WIlnljpvvWfTNVnMCbi03uNyPTdThtxjyoF3ktwN
ViOkuZPBTkaQF4daZTRHBijQ1wgsMz4Kaceail7H3e6ckVssbrhb3kYMIQPrBHDmIyTfAPgu+zZ7
Ell/S/hbWBUI/n8AmR06vacpf+8rZurkLYEAByjLZ2ULMjTvEgieNAXfGrIIKJwFzaoW3EoO16f3
m3fUdZttdrQGmWiTp5dMhEETk8wbtbONb47DNq/myrYejfdJACnsuy5ewiW2kOha1IqDIkQKALSJ
gOVKql5EfEMLQAtdF1DvtytvREKF860wb+d1xHtv5BmRD5dM/OPcSRm6Tqx2JKzQYDLM7BmeEjly
R0QR4z8DCE/21UZ1HmFzS+gWs3HfSZm3SDkcWrcnX56PS6vWnTM83QK2ioq3Z1Un6LgMx9JpMvna
tDGR7AcDD35iH1Kf0mos1a8Gq4FCUU6v24LIHkuuDThz1H48xZetEvfhuo5sUKrxV6xZMB8ppkjH
tGN2tNYG8wVRj5G85OuQEir7TwXw9oprCw3aHi23acTUjYUSgCfWBs8QKfScJjApanxRhiyP4eyu
/330/n75MLsvpArpjjaf5of+EjlJcl/DuR4cGBrvAm+HZpdP+cVEB6rpVUbahPvc2jjgImbRkra9
22IcZEYXI+Lz1vHE6YRhZCb2hZnFsdpZCAVeA8lXbtuIwtbIaBWug6XU0zoeXvtdsTbkC4i+Mp4l
7kRLiZZM/2xeWIrXjW7U8OwfzRLIU1jMo4JE58H2hOr4AFpGWf209SBlIhGqPbaVJtFzu4j/b83O
zxPjE4u9ZPm6aKtx4Bf7YxuGPIGPCq2TICGfuHBCoE8B4sJETH1/J+TtcG3nhKbIgXf6rhI/QqYW
BEfsXoTetgKUAQZrCoua49oHnUc8O5b7cVCjQNUCsjAS15iE2F+2Tm70ijabVRfE1lQqQKFey++V
gxHfkawNyHlwxdRYIkp530opxqCR8QhSoIVsQXW8f+s23iStxKumFSn4RoycbqBxALwhMo/RoXgq
JYELC750xkegfd6t1P1rg7QpWfHeuu2gcm256/K6jTwvX8IYGXkThkJ/KhGQxw2+8W5qpwqRERtw
+0BfcqmyYEoeHcsnJ7MVVoYBHu+zAsJxDj6BWTIdq56zj5fAtblXD94zRgjis/HyoCw8f9k98nG4
h+YIj0VAf1uV77aIC01vLBQM9AI/FZ0aiueh6ahJiL4YZMhFFIQ4fFAcuNanMdXQZviQZ9i0Oygr
0T8EqBwEGB5rGo9X0wdiFWOLq1CSkp2tSfoMQ7/ZLo2sIWymT3atKfWz8eJiQT0p9eKlQHuT9kmB
LsspWuhNsP1bokDJj6r/MUBRpwdlMvUAqlcsa1ZBOnH7ckIr5VTf6Co2owrubSUAcBkLU52qABRK
h9Ep0RzOliibz50JhemCfQ2aEBPBXBW9ky3qhvkqI9rGV8KVe3KaffskYeEHMMbfu6giMlUzJSc4
9NkGxj7Hd5jjwKPOCQrjuiGVcg2RyCc63uU7bbgen7chHgG/NRgYUbDq/x8RaJ1Ec760b6gwnwBK
LLtWcnaBY931k956bNRbjaSV8uDbSo5VYwZaf05lBjbsksBjC5lPZqDGXKJ5Nhqn4XMM8t8aX64v
KfAtVfz0vTMHBbiujqZLynLjffKZOIHc7mlWzNwZMiPkwSDZrPNn5EFGsfI1O6t55lhwJy4oX/Fx
e4bsmSL0EIk2OXDjv//2vVUHUgAvJVDTg12NkQfSS0rRoLahTARv31V2gPNZYtUzpgL9NOhG65sD
+83QlMWTZlqM2OAhzWKOhSAVBoyZzo67YeJvcVxwHcrmI5zt9zBEyUTEQSlxYwSz+lcRrnerOrjp
NIh6Gi5NcLNZvizrlRFYAicEwpBeL3daQXutcYe78TGfIzZ67Pz+1pDMs60vOwu4v3LoDcG9/GAh
GO1AJPCHITpmj+2IirxZBmkYfGlC1faxSPsfARMI8TZ3HYGqpJv1zW9Osdte0N+LXjwUTmGEuL7Q
074T6QJSfk3xdmR+qpr6rAzSY6d5Lx1zzB2NuA9uFD788lnizg4DsmHwXIrSyfVZmuouMdRf/vdA
KyVnTCY3i2DOSLcosqMiI6+YnDzBFct9YXWJl3kjFyx3Te+aqYz50OH5Yrd0cH9MNXTAgdTDzYiH
lEyzUIWp2VGCXnkP7mGuJ8Kw85QSYjXKQQwVPhgNDn2QMlag5JVyC0+eX2JU4LGD4z9DmHQlfshO
pfW6q/DDAED9Tfi8PTWnN6OFYh5eZREt/jv6vSrzvHaQCuRTH6fgc1KVF2TspgH1bnSSlvP4KrtN
6C2O2hO+rdeDgRMcN4Ui9ym840EOIOqI1CZpZ+ckByFfW6JsgHHxYrxTryayHziNLq5h2Ks+Oei5
lWcHQ8eydV/eUMjtGjZ5OIdCGiuZcpMUZrtfA+dIWMGVKoED4dYAVlAMUgPWIQ+QinCpf14EwWCG
waOqSdCv+8hav+UcI8g+/IV4dHJGK353QKW7U8nSINwbOVuY0U1pNmT3L3cEZbwTTJ388/300VWa
hSPfXX3VPn50444o119A8dsMFc2gkJ+xVFhO2HVxAyVltoeXTvZcLo/r4fZfzr5v69gYnPwhUqM0
OrDKGwXcrsNXNttBgBzsk9Qb2nVD3XgKcdeRraoey3op4JG2p3pYjw1ilT97L7qfYy8S0FK7s0G4
kgRLiYss7AwM6aQV1u9Hlg+swO8JxCDf5YoMxJycVWm0o+qNMYvpTKSnUGXlcwA3mOIz3ROhGOpK
uVi5uDGpDM4EfGd5x9riBSHDcCfoTfy7kxlxLG5RH3mzqFClOH8QaUmv+2TvRF3lUXMD/8Lds70i
TSyon2i1PQ4XJX9j2ANOYnUtpc1Z+WH/K0hdRj2ZDBJMmAr1km+B4EMjJ2OBBMTmZHivciscXrMU
JrZVQqpZ/OcFcnGA03RsrcUhSnPmUSkgpJ+4WzUFfVeOwi/Rd0SGzO3+RcGfaKM0Hj44FD8ETPH+
+Lg1mdiIm5PRPAWQilK0lpRvCacyA+GCEvR+NG3PMkWIm9yrY/pUVRD3cOy9hERfyDpcFTBkg4BX
hXEwfLLJuduF+kDoVTE8lqWIQRXhhg4YW7Epjsmwp5lEhMHK0vNYSpAmF+ScHFoYFIAjh3qlqdvX
fLFAdQ6rzNhhX/6lZH3/LAefWJtyyFX6mf0+72Re/J5BseK4rzVksepZqUs3Zy7mPLZ6wBF5mL/k
6u+htehdF+od6EEATDMKnksYgDcYfEK1fjwRJvy8NxZ7kfjHHK1GHzYefQSDUKCj03t8FTBOs7Fi
u3UBKi3OB+v9zbCXwwdKG7HWDLbjcpPVLEyHF7GIZqUcSE9Cc0MB5k5xVQY5ihJulQRo80Qr3AGj
gYuqhYFi/kQsG/lM3jLtEVS5Eo498x+JziwsaJ+ACd+QreNaUiPGpsKPzcC/8JEvBjJytSlDGkpa
jm/viOpPOlruBFZU1hES3bNeDedqaUn1xJXsyfmWfozrzONa6hwcfPeQzWirQPmxKJ+gtYS3lBbK
kXYxZ3GK++0NOKUFywr0c8/HQlOBpmWqQ2JOO8q71Cypv7hKMkIBaIj6HsRR+C1v6Kv6v6B90W9N
p7lttyR8gz2tyCw9owhKEfbbsJkNhQRJ1+Srb4TG0BXnf8nMpcclC+znaQZJQ7wMr4kF2XbxMK24
L9TZyn6klNrAK4XLwN8HT9hKDctPq5BaE94M9hVLP/TEbpZobtAQjKYpuI6FjmMh1xS5hKT17Xfk
m9r913ISH2od16JKcPb3EK8L0VBCcVoaB41vVTLRkZ8Cpex5RisxpbfWRqSBp269gs/tliPbMXZE
cGnFVwebKVJ1pxOCtUdmuTiQLEscjphAvZ1lUxll+/lcFd9bAAipDLqD7k1GB08p5Nhnc7B5utys
V0By/5hh15swlVawPwrQsutfMuwsaU48RRT3fauHHFph9gF+TDsfjIvr0enqib2NUeaexpZngpsZ
2ZxzMyyXu5fUXesNj473q2WkXPJY8aDNIUvJnfzrJ/5/LD3GftcLePeL1UXdGHeJqis1LKPxusgQ
jxIz+jYXl7gBGp5ZD8SZVI5YSTGujSYZA5qZXc4d9DxRKlLcixjv+KJWxWP0TxTZ1JX7+y9Y9ncZ
5SIQCkxBJsgdOVXNjF3jrImGwUXvEcMmf0+qdugP70DZaRb/XxDDyC5OcZIrUOq7frIGka77lLKm
p8QTK4/EfKA7RIWtTs+l4/aILksEzsjvDfAak8WVria+qqnr1XnMRV5hjS0nam1n/SPj+HBGrOep
P5mB/AJ1u7yFQEpiaU0CNsDoncsiEwhauIAIv8eb9FXOAlQ61/tyND8VUylwrGb++XaDiuhWvBBL
FR3OXaje9t7OmJYRdk+yMR8EKSjrzp0LGbGejX7bFcdDYXrJ66LA75FH6eK/u1KaN20psZ6EyaHa
jODQSZKyrpo9sIPPQFFQ1K7HxsQt3mTCZ2/nrahQGD4KLJJNdt8MSE3R2i6Nkj7GLFyQeJxdWTnE
VR2cLNClS4XJJ3owYP7vc2nSafYof8JqhGvybAWC29MsG5sr1y1WAxxelUk6WNkg2vV9KVBV/i4H
p2adAaJKpGRF8C92jHXm4jEgt3OrtOxwwdP+fLuP2RlvbfJnq7wefhQQXE3Fm0QZnGcSWyA9HoKh
OVDvaK7C/zKnwwrbJIS4NLtdTNWrMyQdbcc+CES0lG/X5ft7ccf2pUmBhesVaYpSIX9uVkEAAp7m
x3yQ91n5b0kTujKsONGjlllxrHUrDFJd/SjRHhhJSpLJn9/IKplGbc6Un97YuEkT6bLNEwsgOlvF
QxbRoY6WjyVGSfx9jUeI9iRveSV/ROdAokV0oU2vQiiLLhvHXsBPwf5085+EngT3FfnQKHtsM3ex
KCzWaCha9SV2uxhGr+iEiW2RXmbt94uC5j9pukKrvW81MTAwOebmEpGQSXfFk/gFy6XXz8qyHR0A
7/G6vejzlDfKAFqQdmD3RVCsWsDMHRIJcUD7cjyDiN+9Y2nUCWkq6HlH2fJeavtiu+ty8Xt//TLi
uY0LeSlVAm4GJCmjJ8scU2Dwe/cKQkkvo1alMXWFjIRHOqgBxDFcAhUj5ZQmRe5BuTopGj8UHyhm
m1Kqzh8uLZeMJnm7KwXtv1rtcC+/SpmkIN4nBJ0ziRTA3DtWKZHAGVYntWvdjLcJJwpljiOLtsOa
R8ZS/d9c8ABQNNMzj5BXzyvn3OUZVpMy42PRZWyusN3OEMvXNZN1azWtlOWZyWszFKr8pe9qZsVp
dwm0k6qyWkAil7+NHqJBQ/FttKA344R389+7WqW5bwEHgoG6GBFNn8gPddN7mXU7ghWBdySP160J
gxasACTJJcn9MSlrm17HohAUdBhto2Yb6mJQwD95myQVdXVrDBshYUKwpsoOMsLS/cJw+RFQachK
ZNm5yRP5ND/Zuwu0EGVU01dQ3jI3rg2KYMvN8RPLn+TEGCXbv0FbynDMARcQqzQ8LRjB8PRH0q/f
KiVTRM5StuSRz0YUwsntLPcclBzI/uFZF/WjML19GbiwPQ+Uxv2Qh4xgGxtKP4P2cNWT5r25DY1X
9JJxKBkqTKNQCa/bcwj0iAhxEThcSycuKWBsNH5IqwrATBjGQmEnLJmUNbeNPKaPnMZq/Fc8i27h
yiMNfcBfGPk2Gzm+riv8056oakki33+R3YxIDybNYotaE4SN65Z4avuHAr8Ay4Jg/fUtkoCN8rRu
zf0H7Q5NbFm9/euCVncQYh5S2mG91tibXSkzdsKqkN8LtcylpSXHzIlwH4o33tbYdq/ecbWbioPv
7t2eGmdRnOmNA1nHstgO4u2LeH/nF+pEHyQaD5zBAPNc0Lzv8PiE8FGfJleF5UnrXgjnXdAj6pS5
VT8QMxYjb4az4njSQWj/bLSJcZha/cqB7iBmtf8n4G7Iuc99uj1lk5b1sTn6WLcwhZJQYdmRDCH2
5Q8E3GeTCgYZl3E+56Ee7oBtuLG83SQI5Xo/jTmICOGz/xnjKmGJT5+0NRi+swShvIVDWbmK72nH
LjnxMEuxRzpZsp7JYtcWMYtpbyu1jvGUec6EbM+6D6qD7kuxSqye7Sy94v+NSIaQffn6wn4yz2Yw
csBEmLu8Ou3zjf4P6qQaGt+VBOyI5iyMNv4YnZXBRuhvfAI+9rZjmKZ5a+xV7alHCjz6sY9816//
CpsK7MXmm/cGqkv0d6rihTkb06KG78Dn5UIsLIqAUBIY5tgfH1N74d9AeBpNKxTKh18ZAuFzwYnH
Ich13KzIn7ewFfskGBCbr+mpcUcW0VsRTh5sDyLNcS2FndenoJwdHd8KO8rJFmOcZoMDyQ57fNjC
wUpdG7WWjzs1pmF8l4woV4iHmK/XuWT4qIPOrcNqagso0EvEpM/m4lGlk8K6pzG93FEIkBZZ1Hx1
0bZevvwWImZsSHBeXe8Htzd73dPeAj3nuufjN7Uu7HkXiX2JlulVozxKQZps3Ttqw0gau5nGMDHq
RgA5kgbQk3ADGUN5SXZJu3xusBRfgHwyQGGOG/ciUH/lBuxN7X8LFO6UmHnNTIhpc03eJQ0Jz7cf
+W5BtlfyzQXmRb2gfnM6n0FYc3QbimYEB6nfVymkzuVlTZsAdLdfqAOBcTzixuSNQJEGCvGhoulz
adPxcWIkTBlSFM34lF+Sg9BQNZsdmoCCrLhCtRVXK87N8O5cwHxG2zQRxwzQFkgx0EG66GlzFAmx
qwx47d9CSDWqskmsD8ITtmaUb9i3NSnopzV8TUcU45pkwqnyJY0Ia2Oq0pS+nWRJ0HVk67NrdGUL
nVmnuRCxgoQ4THNvicIZUVpLpFhpDXgTf+yBJ4erbfJ61u9hCYcC72xOponsJjlPtke+pNKkQytC
xBB/q08bCYLLFQClDTEevuBQV080LMkQvWplF6NfljrY0/j4LPBGxKQXPt8Fzx9mgt6cs2/R4aIF
cUAjMSn4FdSleMb+bF53Et9tfUYBQ3rZkyQx9uqK/PgDcAJ6qo2nqBV+k53LJ9NgCHNlnicZAuSn
cPr7/g66IpqNUDH1twEG7jlKssnGPVlUa8MAnqlJTD68phsQqum1XGIZCjdyb2sDzoHXCwdyxJ7t
yy3MiaUoCHOrevlh1kUa37XXcPRAP2iUkJ7QCiOP7odgPaCzgvopCE1NLl4o5+RT9bKdBaDaM/dt
B6tHus3YjjdskOXyVGk3+ZvVW1H5IFoLbLTgi9WvmsoiXPRhExs911ZedUDTU2dsbG3Ldl7B5iHk
GnswJWu35jSwuyZtuQhGWVtymcQJ3cO8+RNl/V9YK1bJNCh61ooYnJOhw4YbIBzKrqBUQnGwMdXS
dxOj3+NP35o2WvCkdo7sSMUXQAy4GWyPbs9r5k4liA2JAQEjlzXncxuXHpvS+Ybjomf7s8ybCN7s
6AsgCvMMaSNmCg0sFnMU2TGxTf+qDwuRl90Ex2kLO4oEz1LmX/hiOTD+Tu4mLR96SKKj5YYBrBaG
D5DdOnN6/n+219ovfqUKubJpItzU32PpSEBsZh4PCdRTo83WlXyWayh7WkKh91c1GGyyG2/8qU6e
Jec2mDuJXQ9KJdcCTqBarp36Vli9cXKa2rXD7oYoW0Qz8R29X71bw3Ytv3EXTrdtg9IorC8KpcE9
nAE15yWOvSeNT9xSu6etWYYKWzP2FjEM+nZdaOJLCJJ/3Z/19qWfPu1+gB1jczU4BNxZkdfC5eRn
JijEuj90MAYvMNM6yjrx+WyAvY2xrM85rw0ceIvJkF1+dgpRVjmnjZdt0ftnCJ2MhSAJTftuI9QP
rvCsFbCKJVH1yEl7odba+Lz8PVnR4T4aO93LjaIA5+jG5H5mn/HyUb/dgq4YcF17ESJHJUGflQQs
o2IF3GIsO6RRUTIl+x/mpDwxSvU1uL6LASH5YEvKBjgKefz/OYOOMZ5HIjaLCMSA+WXiprH7jZsp
fl1UlhbJG7guakXVvl13JAJzXzC0h3SHFQCps3GPEQrXwFzLxKvMLUgrbZPxfs+DKcmoM3+ibIsH
5yXxAlKzGJ42ocyiDBXikmzSZIlN+I26o3NDrj3mkyOC6QSDCQmDS1koiBvj+cnUi/GHwyWGYKp3
HYFGmglTFfNFJj3FAJm5D+J4+QpIIXluiySxJJxtoTyBJ2BX/ZYb87L51NPIW9WDCWAEc5qZQyrP
hpnnYe2Yg0xTVByJ9CsOMkVj+eMsA31KvOTbw5jPjfOaZuCy+9bB/nhNXBcyS7hMc7cfiacsOKen
UQNSj34s9l5YV12eBcZkRr5DoXhmwFUhoS+WDIgbrDLnwUCAxZlCZ4fHzZLkeLDzPhy3yxYR26Hk
ApK+EJq1e5BgaeyVYpN41WCkhBFMwwBj9ROKPgI6Jw7EUAt+9CK/iVe07cNIh2IbxcUCGGzFRnTU
knU3hFGhcuiO1d+nFokrZ34yRsPNCrHqNCR1rYUsiTfXNuME2e8ykMmTbsG/eUFjwBJ6DEah2Ac+
rmeimYADx5rxPDlD0Yp7R0VAssZSiYQ/3J8dOXWBtOE7VZZGWPMvD/A+n39R+SU3mH+WXDmHBW7Q
yxqMr1lFGely9kYnQVveaoEPyROd2nAjuna1M5RHCw7tq+rzc8FOQzyXXlanYSElyMHo2MoXjnAd
ZfTDF/378yPvce2XCirJNsDEQYQiqsDR52RE+/PZFowjNeu8OHyAy1msWzLbfTGL+aYB6Pul0KC/
v5MjSpkQzyeiaV/pFiTxY2wY+uCK7B84SCjBqgbX+nLb+BqLrkSU5eoT7/zvFz1dcEhgX3Y0Zp74
RvwOBdiXqfRsNG6dd6fouHrlx55yxeXowF7JkkuNQ045Ow32ALLjPryvXqNq9QGANo1PxHCtLCWK
AcGWXN95DJ+XBoY6Vu/oKVRaZfi4WFGEkqEKTQWJPnWDqiXBYMmUt9fwU00uhbryx7sHVPawMrgG
j9SLegLs6Pln3S8x1kZ5FKGrAvz4iuNKCneJ/dVYgNYJBZCU3BscI21c9UFIr99K4ia/J4b9fwQc
boY3K6LlFRmQxmejQMHZBZ/fER8yZz82y7Q5rZi8rVNnEcv4LqfoyU28tdnJ8VRZH3OpCjlP6IXu
qy6n3t414QHpYj4tqdwG8GYWj8IV7xndP7yNbfwxhskn2IJ/jO7TSINXqdlIVKuNz4GIamznH6jA
Favx8CDfq0ym2YYAcX/Q01WsvJwbxA4Gscrz/HmNcKMPYp8PTcH4hJKLi28mJjifxE8mp2EsjtrU
ha7npg7NZ7DRiYIP67G1c2e6HrF29ynUnHrkAmXUoXiXnHiP8G9WBUNyrlMoaOObBKy2CY07SABx
bWJn6LU2OK9MH+4BCR2HZYAyUJywru7rnlZFpvjbQTc2w387k1LGid+8dqoX+0e9fH4ZiPKXhoMc
wJUFfDrf8Iq5Oh8Lbig7Z+L5ygy6dBexuM6RDDOefhW8Oe8t2G1B+S4bQKDHqB6nbRipQH3B5sYF
m0Y712h0vEhzPfmZyhPkjQRQyOvjzhDLO3It6H0aHdNGVkg2z4L4pUxAEqoq7aReyBZyym9X//1j
rJATvz40cS0x581BnRsPItHZ0TTBzsC5WN7cGoo3iiyfldTvO2m7kZMIMQnfixQfF9brXWPINwwI
RMaASWCQ+91mj41G8sYdDIQJgdTUOHG1CPCpO7ND0f/R4hhZ5K0jqJbbBlnJSmRKF8yg2vZ23ZMS
fnsidXDxUta3ABCEHLBZHQVdyGjnkku7ydy9qq8EmPuHLwWWapEmSvvPeqf36sER7le/t8Sf3aZV
UzCRU874l1Tn79JK49WMxYVjTH3X3n+6wSXHKTGI8YYjdX/li614owQtL9WpvdqC86PyCL2dzJSV
fVGASYPZdsoM1/Nn2dk2uiC8k9l4j0SPoeS4foSuTYUmURkQqDul8NP+HOm+d1YSgxxpxOHuVQbi
TAQrMInfawCCe0y/Pzr0T37HfLrwDaD2MngQw3qjRT7CKOqQS+P9eenf6kVon/4XdHN+TO9N4XlU
+sHHDO53+rcUppMfMJScYLyflJWeIHIg8S6+3F3nK8l5j0r7LOFVef3jDU4Zow5aVskBJCw+scXv
wZfAGa7JwL7uBgdS9y68P81OzNwkCrhAkGb4O9GmWYNP3/RoVapqCUX05YNYX1PcNH5T4+Y7MKg5
1PEvfkhFBedNq+MnB3AwmMVJYD18715qVPUFZRHXmaQmXpzbypMHGTK9iLq6cgeUSXnmjLtvC6Lj
JjpxCagduN0+UtXQNryLY5sgRE0yAol5W99+0B08tHVR0JoxU0XHDd+JGI2uTfLN7Xu7G6CrF39L
OzoQvqw08UpHoN88ttAb0VzVN8cRZQPPVqa+j7oaRGme0caIDXDADLxeRYIYS1oAMs5fjSdRcVgF
0HblgeGOIG2wHKR4LAMClmRQDZ4wMS+ND+y0g77WMEAX8SnuyQfxmmS53dSuYeAN9TWIulij+A66
glCVX0kHE/zzTtDrm9aNRbrgZNCxV41CNLEZ2dJlGj5237+MhEWZ+BQJfiMi7L35aZUyqhBdAfrM
5t16WISNGeY9mm6uJiZQbBhy0UJsLqLg7LD88SFfC0c3P64+9w5MKbvIZdtkV4nkR7MPLBpll6We
B/nVxEEXMZfmImrn+Y6oRWO68lt/ThjzOXEnl7oyLY3/MzKi/pjF/Yha9ScbNAiHGwN6CsHVJxDE
7mQyJ+jVuvI3FNR7xZlrFTHeQatO0TBdZ99v5hmxvALyIJoUzBghGe50eoRQhpIQJScCRiQOY3NO
Ogd2qxyHAEmbqmHrBgIwsb8FZO/veHa0Qo6iudLC25BK1Xb68azV9Y0s3U1OLwXO8gsZUTejZQhI
3Uy6S7aBzLhfeFvAOJ/Yb9eC2747tbhYhZpEsEYVfwr5N2yN8zEccC0HVjUEOV0KnUvf3f9h3qBv
9SiCpNyxqd+ASQMpwCJIRtv6aL1f9VHYYx9UkRRN4CKSkuF1tFf1IjDPCy3aByf/X/cxfObFcUm7
806EK/r0PoWtQ2Hq4E2CwWukl1BMbKlvG9E2QsaAoBUFkTFR1OJmWDW1uubv4a9XaZmcjXUdbts4
WW5o3rwLgtdoJT1zybWiCWFiDubOpamZX46mujZUHqN+Ttr30G4MMMiVEwsjzQEuNQAQaLc3rDbJ
jaKM//jM8WtiCHCIov0W7r5G+1Diqndej8UADuvhaUs9hELk45V5qNKS/Eo1vml98SnAkWGG7JVh
7CpwONKu9fdk2FMsqj4XHiGxV9eUyYdPYOohVUbhED7a+GSQnTmaJi7gWeYLux+a7k793UNaepic
upSdTIQEeTczF29VSpfobybgEDXtStj+w4O285xWi/zvPnqmf2qa69WAKHXegVifwjAKPbHdg545
onb7T5mZPqu94uOE0HS+kq0fnKy1MlqngOvwK8NehQBQ2MwtOw25VgYxT+C8Bi0YoM3EHljEn4tj
n34zflBu6wokIc1l+93iJQgUQSZR2Ey7N0xbFnED/gEyGspyaHlbSG8ouy/DzVoF0mM9ezqUSgX4
QEgtlXFUnfAw/UjQZQKtRfW7agZyT6RZKkFsgAyBar5jvq4J5FklxQeB5yzpLsHnOQGv/PWjK3Fl
3KFfTJqK5O1qRxDhr/IDdhbM75groteWDj0Ij/ELc67hqNVr077rapMfR0Yt7j8E2TQw8Ml3ewp8
stv7T2Iuogk8g21Z8LhYUr/l7IxidTkecbphJckbf7/eNZHw2D3mWbCGe4BoRxBg+MNFVxoNBev+
5M5NKU1FS5sXO/Rqd+oDzQ5NlXXnmDr8zcRvfo4fTUCVkWeMxqzV9Djs3uEPSpa6W+A//LyeK0Ea
zTPfBuAhiFkIZ5qlRVcZtVpJVlLLK8Uu05stk/8oyLlrkorhnKu+WngjOGEK0ZzZsKXiJBx2YMkf
RHDVsycNuaAW3DbANdzmNU55cWrJhxza4oP0MmbLJYdzhwyabAKuuH+/NaQ3KluVREzsv2yB5NDI
AGyprpQSomcrmB4OTnNFQV9+rQKHOqRa9cCaJ/cKuXxtgPrgBUlffVRPI8K01KypfVLk+haobrrw
z7mvjzTYx1jaZLhmSmq13vd737wR0ocWbbqkpUNembSamJ7lMp4aacgu4AXv4DsQv+u1IGfVNn71
Tm82l4yhCk7S7JOGfBg2YWwq5pd/ihC9F3zsmIIiz1LonwmVSaAPLEXtOcEm2uikYBsSqZd6ixnO
YP2c0c6gMV+WxUWT9BK3fWnm1mXIVXgus9d2rQkIXxrC13vycTf+YC30aLDDCYU3Dm8vS/hKPTaY
Fy332KBQ1aYEamsa+vcdUNgLD3sar3gX49ZcUebGSlZC3bpIGxbZyem+IFZCO6YWoV/MkhvTUR4t
V+7q/iBoPzH9yD5yq4+a8VZ0LDaQZIa4K8p0UfOmBCJDG7dnww0TAJTqQR7Yb7Pi7vvA/my773LW
9p9+czfbZStO5xodL09Y1XjzBpaXTqStzRF3KqkCPqBGKC4cvwXpOB3HlgHQWU19k6p1cx18NUZe
sDdxRRJnsYV15LfmVZvFWDvCmOITpggODqCV8x9OPL8p6N1YNI095LI3WyVLqfshwyKRuV7JenIW
b+WUS3OdcEq0E7fg8NnKg8TnbjKFfe8PJGmo26Pocrf01SSUu9w/s1icn9hwULC+2NBScXC/UGUD
DOrQy+Nkk2bcJxutkTSMyDQZ+rOB1U0+plq0rlQzHABXXKwcE7LzLCCzryYxJTyqBqiksFVmXLyT
aAI0fKtlWNXO7aaoHNvvbOOexVOofKL4XlDV4b2hauRlNVNZO5LOl+q2lj1dxvwJ0epEHjB4kYY+
Zyw1ci61iB8esK5GYwLAzd08B2r74xJKv0AslopBNDheqq6LP+FpgIiDXlQbELTHzsaC+N+GFOa2
IrypR7INdkxlNBXWFjJnzoURFhcpdceuDV6EWXlwysqTL2MCLzLe9GcWBmwmCBocQU8biNscJvPf
IUcJrXfbUTE12cfX0RxtrHoEhtckB6Yh1zJVS848jlxe/sQokfJ9Om84zW4qeeTo5yr7kPxnM5jM
C4F7sFe3XLh1KJHv3FyLKWrelskVr7q8D/TPxYUPXHWK59U6ReIFa9Nd5oHgUhhgqw4V68oVPuwI
vPgF1slpirBIW4RjvRsKbx3OtujT75JS4INPwOkxmXNHeY/K6xnhpNGrzZH/5t3xWgTvSF1ROHYj
QuwqXobIsMDC9EZDx06mySLiMJT310G+K4EkP75QjjN+2+GR0YGnaX1jvntWoj8DctcTgQqM3D65
/vmRChB7/uV7Z/tZYAh6XVDOytTuqTCb6iVhKjEHUBpWPcIorsoYBeIvwLm20c9Od12HxxkhQrx/
m+2wj9UeIbaSNtuNZhPdts0l057kP4dX5DfgQJrlwoVn24HjFzbAnq6g475cBg5vo4PLEVH1FHi3
Tga7E8pqcNwD0CiXBM6mF4MKvmFlNLKtM7gr4i7Zyz23pm2Fz9/dcYcwmQIdJQHzqCsBEVnZgSUs
qfSw7iPdJKDXvmGGnUrQnLPoa9KT1lqT45xfIv5k04rD5+Je/itEUy+Khq8Yp1FGyzdvA7OxUVNM
TVJP2z1FYJgQnLUv5/LSF+QZEelXcnSSvyXACtGvHB0VeSvUPbpcqPNzUhfs0Y5Lj33fVFv6oz7P
es8mugMdUpNluFjooCb3rA26Kc5iM8Ng4JfaV49Vyu3nJMYPpeaUI1dGOCx+CvHVPrxgqgogNaTW
vSDITZL5d+4c39Zlnx/kHQOM8HJGomoTh7zscBz1KWIlqDJrQRm+gETTFAdWX+eAok5bU9QjN1gq
8WAZHcnwQzgMf731GCSGD4nzTZKX5eGI9YMnSqj5k4jHVMuDaTTH9zo9AbTIJexQpEWaq1mJF7DT
+ODDPiT6EansUj9L/JcfchjrH0miTBSgAcr60cIO926PmAWrTJJqAu0b8+Y51QsNOepngXth+qe5
N7/Q+YCxGVI0gRZE1lgPupkl9JP1WWVxcpQPbgN1PyEXCviZUyEVGNDxU37PsCIse7uqrCLSYEXb
SxJfHBcpToSFNbLbnwOTPPPKbz9Am2WfpIaqgFyaO/tGV5KSDKQSaYJ2uFMJOnB+ewzZxS5BoSCe
4oAK/YXkiR5Y2PcI7t7aTEkX3R5Z+xKuh9VqkYLcjjkjrqwmgcnsCtwC4Rcp/t5nqYbqxlNvf2Fp
1pg95U9tOXpR+A14E6HbsHduBz8jQmfpuWy2Q4ksCthqqESoCiWfIkUZUuMuvKPfEI1Gs1PRyyY6
nOrrUNiavnDeS8X/1/M8oXmM+uOw31kJaJEWr2+XuuybwbWkNFHc/rsnORi95Css8MeMvsrummhz
GhVvCTvHq6FNQUSEVgxoIBVYOWilLapMnZiP8UJvKEIMZedlnw8+nrf9R9QPfXuoGDaT2fQe5RJD
986LcHMct0zIYOY+PrRathN/yB9nunA0e3w1vQN5Ri6q7tv7npUaGZnnwVPctLaZeiZcTZz6p7Xk
EZ2bX3upCYdLWcxklQkqdysPdZ3T8CPVYD9v4VzGlr5V+UXBMKCpgPFW466Hdz32UUFhltUlzyqh
zl2EVjNzk+opSIFt0pVdIut5bDuko6bsRikw6f6dGSuIeyuDvOq5CP/lF4Z4Bm1fhE39L3FB/frb
+Jr3DBpdlq6Xc9Hx3h8dvl+fkPkJd+BVlVngVUiAHVL1CdvZthCffwbw8tSG2hH61VY7+Su9QUhv
GuS8nm+mdWUhF8Ehzc0r3Y7RMnL6X1ISPX3QKIUNN9bvtxAuRquuycZiFHKdFvU3haH+WvTXwGBY
0gSvY3jRxxfCjALqIEgm4OjXDqlBS1J4nfxR9jUHxqrnBsUTm9mFtMFY+eoZHQx93OAPwaSeMp+L
cEgdWYIBDn8HUEfsZqdAr77K6+XJ2saHnLpZSBARVa0aM0LmKMjbo4KPTuWNAGBPFfE6kRvXNRYg
kfoOCEuA0IkrR3Z3bcpkCq8ZUJCBH7E2BBpHB5SqIhU8ajR4BIG9+h/8LksglDu9nreP69AcwA1w
w6lUvFyoVopSO49K+p2fm3QMDDyCtMdyD5jHF00U0ZG7TVLwW7wHoP/bOfV1zlVV3LEvvTpzMh4f
fzEjwTSm8KX5IH6hPzzjLxtQpS4mjSak9BJqjSC+ZOHy8O40p2BoZUv1HzUtXyi0o3pLK0YRhbTX
VqFdFG2fxqHsXUl9dtescuA78sgEcAaQpa6KC199DwMfSqsiyoDaTIOL18SKF11pnlS2EE5snRlh
f6Fc2ZXlFVcQ8v3zV+LjVCLdL8gbGuWVXT/9k5uss5kWWFQRVe70apiOM243h01lwOP1P7WcBywn
8PSspCdVCe5b9Bcmn6iLmt3UiQ4mzXM6+0hN89PfCJEzxYXuZbUmv2exTmwD7g8Tm5AB6iexjUCC
gxKO+hffbBJGa1uMTfVJVH8O4sNsPvZ1bMI6lF+FLizBgBhYygiMQ3cFXHtOB4vnOa9Dd7CJLKOG
BVq6d2sZmstCdr30b8WSFIY12u/rllF/6lZ5AE0WyAt1OLDO5HS9AoNszbPFSKrHhCeji4j3CdKU
Kuk6PCRc0WZ3DFErObMa54GCE7C/UiGYRDVuJmu06KA+T2mEl6MWS5HVALE3HXTHrr7Dj0Yxa/a9
Z5WO9oKIF3WL/osF8krbKXWsvlMWxShYgiksAY5KXbyiNl1JLD6muHK4cbUYmAA9N3kQ2BDajwJP
vkMvqQO7qS8gJLuhmtUbTvfoVrQOYYvhya3/ygklAo3uAisAfrCjZtIh/zXk+1IMMzmnJKkRFqhN
46H6kMbZh2V09ITKFd/qRoU//99aVEqTE7E+D6Md95XdLUUlYN4QRoyh0g75lZzGwebciDhQttTx
f+TA38F7Ojs8eszVORc74XN7i6d7XHYWvjIRkgpe4aTJubcXWx8LrRY/MoMImQ7pbtdC0YygQVWi
ypv4IaPvITIfR2o26U4X0fGXQ6onMdl7E/pigu7CCYFtoxaIRX2wC39DC3T4YxP4Yujyo+L4UIf+
IzWVzzElU0echkMME94BobltHcaSJ7Ton9Qa9BajnW0V1ZGa6PPtLtEdMw6lrmMU06LhNkyHToq3
4hRrqtvzrVUqq2jdcS4UHNAUUSEgvMkqFdUGt7OGAs5bjm1xlDtRQiXJ55Kuax2u5qmWIfbeGm9y
OOOekhmgSU/nhDHBRrvNHqSYiJVPX92PsD8OUJFf5RuN4XYOltrAXYXgTV56T9m+kmMFGzuAj/EL
SHvOIrhRtrRI+fV0NU0qM1cGM+ZvAGY5PfpXzFVEbCMwzl0ZNLQNMdENa4eg8cU9tqCymgCKoa8g
2nvzkPewHxVzRS6kzk8B4GCwyES0s2JFd6mVTzM2sDSqpRz+iisZKBb0JMT7sBG1r62B3ARRjY0p
+VMRZHXiMVK9vXCN94vwwG4dQzb70/peA4Q5wxV9T1xiYXL5MvVZ/C6TsuWb1scTbcJrjRLNXcfH
f2jkMH3peVi2DM7iclB6dgBJjmiMrcp2VFXJfzruUIr/2fuB4EHula5hVacWq1wEQ4oh2tNJTLu/
aggcaQ3QZnrE2FcHR+9q1NbZUdWvLcQG63N7fPnB9clTXwWWXVDHBSL+wmQlqXYlPd+F0Y3mFHFo
K9ZwbXJPsU2d0PZ0JmCWvTsYu7A0LfBHOS1YKp/WO4jnhOm7DhktPKfD322AvAjBEj2iozSRMpTc
D6cc9JwQ+8oJ2qEnRucwub0iTXKp3fP+tL+7F1suD8t7/eYyIPier5RB+fGJjDwRG8mdX9VsptPI
rlEY6ok4LGiq3G1xDvXapbNNRRN+LPLA6ZScESKIsIUsdElW1hWQOQomg8fGie9wQLKfXaUYmQzX
LMmpO9ivYBYTvD6DwmF9zIsgvN9rhM//OCKMtbYrDjta9eHjvSmu8shYb0WRgiEBPFQ/sgf5WGAd
4Zw2M2hYf63Uqrh2wgMtKtKw1na4E5JguC+G+TMGjZdbmqiMca7iO24O/wt7gvHpHpwgAL1/Ivq9
0U08RLySPdQgkLpngluaxhhtcEQ0GbtuQfC0RkkerFsXWLt1Duz6783Lqy2Ci2BA6F7b2hZYIGji
ktXJo0FuUoS2eCn6g2/Ved0i8lw1vDkgy9IJAhNzLhKLkqEYmZkqDCK8pAI/Ktx5MFs/9MYbNWGu
vj3WpybxnEThWcuvV3wrx1pGP35u2GS2I3aqJno+dE5TMZP2DHVR635DNuyCNOtgG/TxrC17MGao
2xaO9HryAs4cM1VWn6e9Pc8nLFfkyW/+rU9oodevhaMmT4CFHzePA7ZCchu3aYF3AnDsy7YXccWF
JzbEfury13T3WZa7Lvm3RYSq5hZKSupCmzdvcPDN1ct1Qo26CadzMzy5lfJJoAukRk8WFX7XRqvH
Xxhfac0fWOcgnCe1cVXBQ3z7y7feoEfhs4yWJknmfsKcNiW6SohBIIWxaBxgOK1Q9qaD5TPLPA8b
fN+qzzwDETLc+f0iiczhJJFbcymJlUkXQS1v8S7iMUI3r/a+4UkMwX8jcMenQW6X59Msm8B6f1L5
YLaFiaQhwzK0A9/bXummv3SfNnvl29mHiLzND06ScNZVIm4c44ii1cJVUt63DW5EmT3IpIWsSbck
SNdebUG9oHTNo4mlpe8nKwf18OsPIXcAmrqXeJTilQe/RQg0zDXdB/sX7NhpSu5EZEl+X9OZBm6a
fZ+/pqfK7WA8vQuoILYUHaszHU1wLY+rwOYRzlQqQRv4DOqsT7+AWSAA66QIzOZR3DGuDJ4lzV5m
p6rcr7kuL85pNngRKKIRT0YiGTttgnCtnVHMIqQ0reOcbhCUvHZlUePN2m8TkIvUNMjrOMtpfKZc
hR7srXZ1SCzz6KAK9MIsGwxUp8ovfmwD3Ko341pxn6LYp04m4HrVJ7zCdQVF3AV0tklAVgthk8Vk
59LA1ymeCD9OmLSG01lchphk9WO3c1ocICGOJtAOcDQPT+YMPv04RTl89Av+lu//uRYor+ZGZvhv
x/e6pjcCrTXPT6xF2bBHDnglQzFItXzplxK5JBIutpx8BftdSoU+hgsOuclTemLTxje5uP1kqGcM
argrdLaHLyZbAI8mcAD8AEmGuP8xicIjrJRPs5cjyHlYn0kXx6XFQQ0IIgcW5q+W5eT0DTuDa1Hy
/Et7YJCqwfpO9ICzXoxIR2PavkIDRQqlAo5TFXU5puEFhP8SLEJm7r/PiVEtQLG+R2vE2Fz5TBi2
AkwJR/SVgmDxn3jYk71htH68KfpeTZ72YdfwSM3OMNrUyXIXnFNNxb7/h5EWnZFbPaM8ef+kEfEG
EHzHHGfktSxPU8Ty9hC1mMPUTrhr+yXsQBbtNFUTUnpw2f0PGp6LNeu58E22sbVqAQtJ1IDte7qt
Ma3hxOrotVHwsnCuDBEtuugzoaTknbiP3SbEbVkTaKj9p4r0r8kMRbrl4jNwUJ+icZdU7LVdicNv
l+NigFtyKl5aAqrjV0PXuhZVebgLQvlmvoH3hbv90b/0Jts8p7KMAQpo3kfsHQtqXtIcQmA+/fNp
2Koj3Ie/rZoLimP/t6IkaWHnI0CyFtXeZ4tyid0dKmamv/qgIGJe7g5zadw//kQ6LeE7XmMAlALm
uGPbh5GayxI8GngFgYDvu1yIYN+x49KJFijoBFzDkQT9sLPgcg8Ol27yGdM4cO7W3Z1y0v7aRTvq
0POtYdb8fPzI1qKC5DCW2FOb0qkq8P7v48PwFjkYHSV8YDSi4qMJcfW1anLB/IPWkIej10Kdnk+O
8wAA1l2H4fpca5w2MCRJSDiuef4K3ScREXbp62IDp+khFhf2cvGDBe7yNK/6JxKbzYcXyDBIpuEA
Mx4ijVYlFzUk8YOpLuMFAWk8R6yPFDtlWY/KiAsGOZ0/Sf22LTQGRFad9jTH9rY+X4WrHQGXZhHW
AivpB5RldDVXiU8WMFsSaYuwZZZokN4JuPTvufrZpK5GUUC5ovVSxxAC9WFjbCKCPl0+29nk4ku2
y/vFDqmRpSYFCwtCMkNhphjzxDVuUL6103bm23098QQ/ay3trVWhOw+gneuWfNafq+9XHDlyacSH
h9zkXGqTpPqSdhwz/4OcWj/CCs1uouL5BrY7yiPkJVz2HZfFzmQq56PZUT+p499c7yb0b8UiXtKw
jx6OhKg6AQapGMk28+cmO7x/HqjGuKBqhK3ngh1nJSwkCQghOHxCjgP9esQBsbIP6NERW/6AzroN
0x86JMgO1zwta0ehGLSe8RMu3d9W20CJoBt3wzFrPvAdZE1UVyE2nBVk2HcUIdR1G07bCRRKTSul
jO5tgEXW73uuE9n/5xlcYvfmKcczA2+Z78xMV44qtprzP5/W4UUWiweSBNQg9oTnrz9nAgC//n/k
mdUaQxk/5PJEI8BG9Sn9SY3QJsiCUpe+RUWuMjM7sNZgycWvcBEk+2xG/iiDzf5yqD3YfqzavE6T
vKlstU8teOpYcR7lePmaEuEe0eitAQpWy+6gyilmWacfIHDhL65PTPityMmVS8k5ShgNl65DcRF+
M/IA2g4hm/U8XgTrmIjCDbxtpKONa3vh4IQPogjx51WJpsFqvhjiwrS1wcsX33N5lEI6e3VDo/Ye
n57wlTST6D22ie3DPWQ/94HnJpDSCkp5XsQnsyY71UexE7Ep4kor9IjH9JfuvtdjZ0GTKFeI8cmJ
L6NJjtaqqS0KNi8X0FL984htpT1wsj+Sl2DVgYbd/38isTDHDpje4AXI53Jqq8TMyjuK1WePopZq
2HUVR/R6YzI3aMZjSsdapoPXSTV89CZlDB/WLj6AuqR1YTxgX7iaPMX4MIWsZneV8spniQ2uX8em
wV2beGDrv/GQVSeD8cggIXfN13dhYrPokF0tNYgwKbNt1QN3Wdq3AG4JUOyN/AFUvNICtLc2sdpE
AOrZJpOpKCfZp3XItoJOhQBywb2JecD8jKebTrIGCy/fdddhnPTMZOqk/F3ZwCdV+A1lxAH/rLy4
1WuPZigmk7l8mLqKpmtcgtoC6eNgLQ8icSYTMWgHwIgKzTzy1X0d7WMW9+wrN6Bn/i55fSnmCfj1
LVVE40NQVucsgLzQ0CIpDHkaecPMp7HrkRxsROySg5E7M2hg/KCsLbONaAoa1Qzz0ehsT7TZUorL
erctGNveBZ3SJANXmwqJYdR9MOim5hiP/FJOfoiD55WjCedyu70SFybgM/c3svwuuGh3Sccs7uEk
PGGD6j3HFpUOD5LJwwWG0eP9kmkncUqrGo/gj3HaLC8bvPLbuvUJnF4y+Ps6uINvItOV4o8q2bIb
EcAfcFkysbT7X0SvDcfvdj7ruGj+KNWBduZrCOebBOYNnGPN813bjDMKfbuPV/svOcFHyjrxIe1V
X6fza3V/5TwcHbp4qhH+EXGdjZCZu5223kca3n6mRJH9okww/UuXe+aZm7SVOaj4LZQNDXeG90Nd
fI0qgL2+b05h1ItzIxHFwwz0ZBB/LlHrVbG6XAyVnbVlkf3E4IjaB+6EaSGCO1A8yhiNVcGNNW5h
asaZunpqPBL4whYQQG5dETZ/EiSe33S7RsrVbCCFZgnOLh6eK1F41k8fVFqnUDzriUBl4i1+aAxA
bCuWVIgVZaHT1WbJbkCADpRfv6wL543DnwoymLF4Nxo7pG4Qv3+EajOalz1W3RzOiVE/St4/NtQN
kyAbHXgQEQJCQ1vXVkXrBYJFBHdZiu6Q0DP4CotYaiV74iX83au7UFZ4kye6gIAMGZVHfUx7zYSB
oG1e6dRwgxgJR+d6XSf81Nesi4y4IPGqc7VXrMm8k8W3NYy6R0deB3BhE6cqI2G6vSb6K+87me3n
6/+cfoUA1oYbj93X+VAcLyWGs+D52X7AWCNnccqparyW4yuTiI7AlpFz+vsVj4Hhoe6UrInaX1yg
TXjpLa/JZ7DlHqsJhziLBaOc78aFhKurOYB73GXFkd2g1OUitDP+jyEfaRg+8pNuhhS+06JlJCKP
A0OHt822T+38QMkXYgazceNjh9Az1BmhnxnMUQTxDmvvN0uWnIPwb4B/KP1Ik6rnlIHmOdXDyPgz
fLhpQDptXzW4hPmBfvwSUeEvdBTIyegpQRm6oyNSr3/ucMzF1o8/ZEOOP1YSf1RrRUd3csxsVezI
DjC2fvt02io4zNFKiZZ97UgE2Z/YVxbo7Fi5xf8Frk1qN0LSkRLaV4v3JQ0Gdu3WRAaQ3QG59I3g
iTaIwGRPfDQhzs8PQprzD17IvssHH+1pnWbXPOfdByiXdCPdnW7PjN97Qxmp+Wlc7+Zyid8CrMJM
jJwiYWlhyiVzYStQfoLN7M2iJiiluDH+6yiowK+ztv80MPihHd7yw8nEOxNBCb0BoIU5xYxm/PCm
JRfSPLiLfL23AwcaGE4e2YJg2gqQwGQyHdFG7ciWnkc3joA29g9nmHqtaGhuh7lLWApgcXPx8uE2
e45qWeRwTNuGBgoM0YOc4jii176oNhiLNUIetnMxrTKuDw0X2xhwGGJ3U+vFm9oojwViE9CT9m7J
z36tT+/oOtuqye3B8kAjgBbeb0upT5i5oHPW8E2pVgSN3sXzdJuhT/8LZLww/ZuaNpGWB9P1mO9s
4psOMfjwppxAiHa8PGkUMGTPqORYj9kTW9IcqIJQIDj9tYBP5br8EsK56B8BvXkLeRsv3weQjVAk
tmN4rOlEbUkYNHJ634VXe6br4d8Hc+M8xtxIlusyK2Mm1bOMzGSq9dBsnOXJaq8+rfzI4nzR//O8
EMhRSGRJsLGI7LTlvejgT3FBopM2/vIpgScjwUNT7G5tCi4d5y8Ua/DFe/hSnw4E6iJra5xp+2Tn
CeXin/nFaJfCxbkoi4jC24S7rfcczZBVJOXFOA8+VCB/sxCnFV1vz7AUsREeF2cHsxiAxF1B4FNW
1ruT1oepeiriV72Ly6313VfNo/v/QvN+cEvJ5pxw/poW8oxMTEtejCV87thkQfQr7ATBFYxg5nE+
1Vid6ZjDX/M0vZJj3nKftq5VVk1qid9k0wNNMY6b/xc8A98WpHUD3yz1sEIgx5lsyVHUgHzH56Pl
4BABtVrGmAyKfVrWY3gywpJvjvMWJMgV+lvY5dtEKxzrA4JNY/OppAS8Dtb96w0X0ROvaSl+peCq
nzdQ59VtQhtuDZVoWdm+YTuR12ofFS5qKqqx7h9K0LMXfd1MbPmAVVx3dHuPcwPaOciB7MVXCc08
/wB6miANkP3Q+QzPaDOU+T6FqrB4Zs4Niz9zN9KE5GINueUy/Vzwd96IlZzKDzAtZMd0JkP5EnlQ
nprAToSrzagz5j4ZYhVgoYJYLzjXcNyM13+l+iWwdXWGV/i361NyDCYiQtGP/i4ZMtaCDDUh7uK0
alAFOg/1VzCZS1n2mZM2pEjLbT0VECNkAeCWroft8I32LyzoHtKa5IUgmW0NaCwYYYmohfcFESTp
w/r/BcLAVkPdyEo/TJp8Gzy978DtDi3/NF4TxJ6HwUdZNFFtRZXDIAnPwk3zA3/5Amz0kDPEaOIK
UcS+yqOdYd9pYeM+iT9/9rjk3SzrKutpInYzbYmnbDMj0Tew2tJU8CKROZtdv/ppwGROfPL9vC/K
WvZFbE1vy1p/E9S0X1GI2Yq7fMyWmCHjBzuojTDfFvVURaOhNUK4rppohZZCWkhAeJpMex7EUwuW
QLhQwXe011JLV9eUoolzx8DxZ3FQ3WjGTBccnmOL/GlzfESVKwaaII50HFDvU2Ifc+vnII6+L5eC
uQDEncYU7uyebvKwj9HAHrQNd+aO5Df48PmOSUiUH8bYuVstDHyyHppF3gRawLJ1FvbQZ3snpSkW
ELzbw0f7GqFqbHoPauSk7dZu1y+PCehbjlJXTGpCtW49oxq+K0aNDWb4+iN5twyw8NA/cphIMqVT
wRWC2yhHBwq+NEqc2qX6mXKVEk7ezfj74DEpRsHOspKA1c9YgoDxr2Rzk8VlQV81OnmH2pbWXLz2
Ivix7k1j9URp6L8YwlTmY4hU9e9dMARJf+gO0Gvoo5FCcFSdJzpmnEevRmqTpiJNpMt8x58xz7um
0E+0/KHpyWlJIJJrWCrJQct1ysYC3CIwm8V9/0NDff5RYVj5ka+7L5/nW5UQuOxATMHMkbgD0YdG
BKD29sc3UzE4EEBCcafC7fidGUV4SunEiX3NyKkgDhyaLTD3FNOZbsYIglI0VpRczNAjlJB8ZBsP
1cMVyW2Nu9dvnnBfmvtNZx0O6b42ausAkjetfs18j2voKgdsnH6DUsXmb3x+04apNV3MHKbbKKku
cXAwQyIfUtAXtZ/STOBKMCYDOngKqq7V/KnpKCt32olBa2S9dSuRQsPAVdO1hq9r+ozZRShutKxz
Lk+GUiMWa/uIdLFjmUJBVq4zFk5altmgcOaEugg4+yo28Fp6xW0aXkuQ6L7tQsSv0ZYNWTUJeQoS
1bJwYVxoaOuSl7OZrCzB1iWLmPud4kec5Y4JA9OsMZetzISPyZRclc+moEcdAo4ElrkJ17eLR/+I
UG8oLtUy/D9pJaY+oTWh1CSD3qgfD+3LbXUrveOta1fG81QAFzA1rT6oWPcsBpgFuWHdZA25qWhm
0fHifNfF5ieNVn2YIDoSXRPoT1VPx4MYwsjizzGZ38QzGNve3h+iIvfs1WXWubPCMJ8qdELUoK7O
UG0tCNCbvo+IJNElzrZHbCuuDLygm0eqPB+tiZRq+m8UiX8Ei0TayjbFSyPzJZfQYpS08PhwkknU
2daU1Zx6neSVAvhtKh3Ob72W/ugB+CzWqXuSC1SvLKOVhYWRlxhci2OB24YWxjqakK8ZUaEqJ7cN
sjpCREi1oT30eTVYIe6NTjRy+Td9r+wm4n6LZKiD5RG9B1H9VNAVZofNpSCMADNJEbqWfNWvljkL
seSgqHjpiS1mNq0GVCwuXFRRy1poKgMAJuc/TosFYVMaCdYM+kFpZ+mvW9NN9C1tqEDryxptsWka
1eJNb7rvcn7opK/ZNHtdgTrUzO+N8nPJfaUOntmV0Q4wzmLbIYYdU9d9koZtLp/BUD8JODQh+43U
csxkLbG4gyS8S04rnHDPSQQgCRuVRJzfyg8YWt3oaoyYRtHpQhEa2sJ3g8DHD/c86LgOXT8qJpA0
wIHDOyX6VAeuSBZpVtcq6Yg8z2fTXELLm5UPx1T9UBqkeo4wOs93019jI1B+SIzEgJ5Khyp7/CTv
xCqtxJPQxid1vlk00Lyx0j1Og3rV2Nx1iDC3LwFgaTu4eRDGmad2cOubNV7HUrH3awnENv5e0ZmT
KXE0SFECWm5TN97dZC0Hwox2LJSFuCSDbRYpLr/TsaxUS5C6uKjhxY7P3WYwfa/2Ouc6xsKShJLv
OEizdqG1RP3J/3Q9XWiwjl4i1uS3sngmeIfuu/+1LSzRrIG6COzd377Fufa/2KWjWpEej3W7+crK
hHS7vzwv9H9mVRcqLWkg5s41XYqYXYUfylNeXF3rthPVfAr8MZEV3/5jkYnBSW1NvIm3ryv/m6Ou
G6Q2sZZGAZxiClA8MYSzYaR6mIDCt8J7ZUqKDDxJIMjtX4fyPN+7pbxMh9hBUo0LAWkab6bd9H86
n9k7KnZsOZgvjRlwGRn/jK7+w5bMKziJpCna6zA8AzBS9WNaEom+8MTs3R42J1Lqp/mHxrWhPr+4
gBp5C4AJAFcXCwQZREGslOBdto4xq7VHizNU9MUpNzw25N1PgDziSIrDz4txChf2nftcjmVXxd6L
NnM9x+mvzoaBNa1PcJpeYAVIrOjKezh+tA+nhGYLGZH3v5LEoXoXKo9FN/WlM8li+Hrcs4saldAA
wKDxsQWryaFjJJjoCsNDJKH2idKeocsB0kIsfIbfibkzSZW93lRwZPoxkZNjMU+MJJokkWC0uT3v
j1It/1FKAO/jeVWzQ9W9TlxRQIn+E+Nj5Vc2VJVm/TMoOLGM0qA7+aU/6w47tOGMgeYIP0LnCGZm
tNIipj5oF2IfNUYN0eKt7mwYvUPfgdQFdb4Zm7xftj0EU1h6MLGjDFQnnmxo00EkxqGnpYOKm91s
EwG/+nsijBP6QmfT25Qs4N/TcGrDwY21lTVhVhbw4j/bavCdevEKcQzTtOgNlVHMgkiN1mvUdh2U
qzHB2kCM1rMbK96fo/+uQwoEgQk0Ymp5OTMAIavpQLaMikaXkA+1WQpTREW/ATvEcTfvXJ/qX8nV
5ys+9qZ8S/1SjerYv8n1qCe0yryC9L3IdZRvA9fqVNTau7mhLvsD1/J0zGni/OKFyJ+Zv5mqCe/7
vYtH7EWma9AxUhcMht3pPXOAOsm8LqekGa8o+VlA4eOr/67WdmAd+2jhiEvLigOYIuEmEYZlRjbE
2YYox2iaOvikncoM1kVhW1VdrabmhYoDfuzWbXeAamPKRHOd3NndY23pajWOuLaDFSHFE6zjP37P
HKzBTIKhFL+2plcBsT4kHaXYBzpT+8SG26UdkqT5Kk6GyL5RrXR3GGqaKCbJott89DNsbfZtu6h6
g1g4IqUCkkQtZT6q3oH3AmNffNlYMB4uNkHZQ+0xLQ2QoegH5RDC3JnzcelEGeb4yAsg1PGW3lRK
zLFFJ5u9opHX/FvLHW13zYbdtb+Tgzrc1FLQ2EJ9bOWHXx/TQlX4Lujg+XZ1CA3uMz2LyX3yDnEY
WKpJ3hyDXbmPHqMdUg20nPOykCC9rswIjG9+GO26zAAmQFgkbunaeOIGVuOm+kU/LzXfoFJWaIim
We3pRva9ntK8HnMVtCP+VylqBM12NgKLk19jZ87Im0qTByxn6ioqeywdtMltx9UBra6eZonsCFF3
pYtF+REDljtx2HZFvlM6soRC+o8UVlAZ2sA7nAuqeRzf922fSrl6Xb+dp2EXdwMZ9c0euRV8Ly+x
N3SlXmc1uFc5pm3FbOk0u/SwbTsYsU1eWW/u4rp7B5V8C7nG5P6RAKSuaVb/rBsBK1y79q7b2jra
MtSudIxErTEWCkJi0dfj6q3lAcVWUyK+m2S3+izByC+LG1ITmSX8X+v2d+tQZkpbhoQUX7JR/CUA
74oJEvfB6sjRWA2qkPYMFBqkm+F41R9uVryjMQY7p/MnKmKh/k5GtflMs+YtyeaK3s8UqkiEzxnC
GkTGCB48Ab2QpLCiPgrsjEBRc2S9+1aV7ZNBzjQHCLYLe4i0QeBa2n8JWEfBxa2jMPsn4DdpFdfS
ZqiPdLNMj+ULrdSpdqhL7lpLT0jrlG4mBXUI7KmnsDnbwHmupr2RwSkPA8VZxUTBo6frFHNKrF53
TU/HeVUEofspShx4D0znwo/BPfjfzTuhGmHv6Pw5NQKCM7+srPyLXTCxBZgUk0mmhRFb1VKHdn7f
vZ6tpHVgETMoXT/7fXjR8GEre49K9Q1FvwRafLnp+f0mQSmE+9FYqqkjlZqMJLx9E3CkpEjN4224
DF3dr9YyXExT/7WwCFEyFdu7TOCkV6oExhkRg8XUFZjbuLihEjwvVwuWtMdc37bYSERIXY55cNa5
Ngch8TGucz91soMYKaV8YIlxMHNaodoHtk1j8WC+ZM233Ni73dLiczLcM3NQs7PJi+JrgOwvVJUS
GAbnlJybAIFRfNcwNEo91om0qO73JY74zcZ7dAAHDsq75T3ndv6S9XZ8tvgUv/mF9cBc3M35rSOs
oUVliJoxyR8dPrzuw87hS6ElIvBt9CBJbipWtGvk0ILgHL21Fplpqh/tS7PBMpxz4+qPBnwUUq0k
ws1LXewt5T7/+d3Q2oLc8S+z3mToJ4dNxWbQQg9OplZ8SnNsZrXXCRrGOM827YEvCNyM+Ketk62p
ezSsOuf4de691SRjjrCJdGvBG0sp5KBLykRKquBBxNU4F8TVttEHhhL+yTRo/OSriY5GiaycRoTq
UNuVi4HSuD0Lp4i2NWkHxZwJ7TpT7XAp9jil9QYzcMNFsaDNLHBlvwokEauQDPEVssldOR6TiUik
vevGyPENvPDlDWkm4rSJWrb8GLDPnHej7fQM05+SzJMXWRqxq+1PWpMNSxuEc2qe3H5bbx8MgkYY
Rm+joh5JXYrK3Hv1Twa8VtsU04FCVJoQtQUGYKAm1s/l8iBjoXsBBvZNoUyzsUEZt4sUBgAcYXVR
duf1LbYhw6/fxep+W44XqfHVuxYKA6KxCc1jmmWkoo7ojneIWo/OxYz1YyRFEgBNlEjUXQ9ItHfZ
zE6cKrDQzd3kfE7DTOU1s9VVcqKtzdOe5AIJUubYflt3Ig3qTmgECTUp6n5beBspGRVsm+x4fjAY
EcEUUkV3xmYRlEqMUm+/KXqtlkgRuvvqlXv8ht80fACftAEwOvZuFei2ui+t50nbNJRLf9CE6Osg
EHhwqR/7N798gKbs66vw8OULC5AokZ3hSH1wtZ10xtCli/dpnz9SHkwEv2JThIDFUAkkoldQh+Pb
n1tNlpwTbPrv4t1OIHsjt8udrlg4GBEtpOuZK4XYPMJHFm66635EcJeSaJ4u/xaflVQUvhUJfsmN
ySDkccBV+A7F4LqKZLsqnLKksd76ikyN04wy20Y+JPD2xZM8vWvxxfzqjz74XuIKTkzSDZNb6GMS
YiajceBHvR8vrfbmHVtUcgRQzPb9/lyU/vt6zBfxM7NkTbPlOKjcI7oHQAHE0VZrsWPMUc0Z5jnT
ojwyXPv3wYWZsYKrd0UdK/K/5moYrZXU2Q69qeBvnfC2S213P7FWr4pQ3sq2zKKcz5w6T0+1Aov+
/t3pP75S+l+Mt/JkIxpGQBdsS0PYw0tFSC1PKGpOOSsztu5HJJGn4EUHM97WPe5izkihm0KPOaP5
Dheeoes0iZJVeBcvetbJBEuniTxyyYAr43tDIl4FmV8kTwAMoLnw7HYLU8NUnLiwahqYcwAEklUO
YWQfRMjFEsrf3umzerCirff8ROrFXK/hoTw0wRjc2v7ac7ssuI021Rn5yB2f+KC3HI1udlH48LEr
qC4PvqLBkkySswBEmqdifGFXsLUAsBU30RBsqC8wOwF/pd8EC3Oj3YKaTUd3XlxZYI3/hyG9pDVG
vrGiKKQXhXHGzz8yx+OYqIdmN4VyjePXSf+CiCLnei/BQXjHLK+7c0OYasx/++GGfw2Fu8FDTRqx
JgNVtK3Vct0EdEZPUwMtG7pMJ1HA1S4bah/HafHXlMkXdXObIWTEQ4JPe7p4yt+VExuou/9KbEGS
/8bfG1JNDWcdsrh5918h4XcJhylUSPkNUEaUFnE+s4D7yejmNj12HrGEQXEfpYV9EBh8wJ4h/tWB
8Wb8h1e0GO8BKpPyN4Wh7xXv/ebToqYJ91zSgvDEOZP+3oO+7C+YySeWahCoEoIIM7zdFyucZpW6
GncyC5qcPfY9FD1ubo34ayDKghFXeMP/TSMFrfD243CU7MKXzDCZtgOpG3V/Yha0X+cDdfwnYrfl
oYqnjNnD0sjt7oWhuOSf4jAO0CiiPtNdkDhEsUEMyIEBow/r1uMnnczOaOo1DKNk/tg52yKY3sFM
tZWgGkFxJx8D6mZbn7AvJOVXDEBf1iIrgm8QO6aln6DIsIdW+lC9hRxBm3K5MuMD+p/kOVCd22Zo
ZWJQQsANF0MdwF6twVXPZ1/e+7fwQjpE+TnQQRnOnf83+jpOkhllo3pRCem+Dk8OIVaBKE9k+c4Q
Q9GEtsSJJ67BS4P7/cqFNahOB8uvHD0CuIBlkwy11ABTK6ULIXPYI4sGFq8KJvBJyd9bVNy/klxC
tvkyYR8qdrlVFz5fXwOJTg90o8dqRVRhF4LqVkkUrQE0tsjjIW4xPk3MXgZMn4I7I727bsEpxLWt
WAXGT55QHwZLqcLuKv7Qpv2PjYRYt59BqPzVtsaHp0OhExQ8+XzSDJsFS5ALrNyDToMHNogNNF6O
HsvRJ518tywrVx2be4ismkpmisX08s0f+vQkhUUCZCrQkKfXEjXsgoTPPQlDmWOQpQmP8UFxcOML
T8tf8kZR5PjGiVjdrm9Zp64CBK6FsOG4A8aXMOsAN/YyiCWR58BFwKnCf3DwE+WwiskNPeS8+Qak
S4E8/Z86JOBWoCODBP827r5i/qz46O70hcJdrp0yU+jvsu0PZ6WSIcOouUX5wwZdnKRCDumk8U7e
yhdtZT6NRBl9KpRa0t2fKQYZWomoVe3UDZqu0yJEkgiCHHVUHioC2tIKE3EEgSvFwz+RHBFVC/3j
hpKiPDx633mWqPuQMUwmdFtwKubHnvVskCAJM5Y77TJOt2SYSXNsXH+icWYFKtIFb+flUcRxGozX
xK7NjHBxshMwT7fW+pHeNeAOcrQYOoTY49l107AszfqFshgtYBY5lKuUIhNLXJIyA1ia78LLsVYt
0694qOznW4NU77GXwIwq1FamqAu8WHoJj6r+vrTZ1yeTbfn2ExyLVmpaFINprUWGXJC5m4/mDldG
QnelgfZ9tnh5hbusJq/N/RjY5yjJDJA2Z5vonBCZ61eo8EWumPjeMwErfhdh9gFPtvxNJlMQuc57
tPsPoj5X6tpgNUj2NsU324fAtp4X3z0ts3IDFqCItGLNcHqWj+LcOPIT1WKoD8i6wv7tFhWajYpr
JBlvGYOU0kaqj1u5Lwl3qASFLh/RNXSIZWlQccjVW5qdz0UMPIOtShndhBhOKIn9XYxZb5gFSaCZ
RVAi42GsIRl2nzTTULzvWoZjVp2G9Bkyy9yCJIyi3fYArnGgxb58g4BplDLtj5jb4dbHtCpu00tU
97d9dk4OlVHJZSTsM5gb2kJmxXc3QDFziLHU7S1M3pLsRPArZL95AX09/yC2i3MRE5CSW4vkYD1d
sq+WCoB+JExhuljzVSnCtw+U2mDYEzJ0lF6UBJ+Bjblg4RjfV6RaoZ0EpeT1md13UzAP5BrP4f3F
eFcpiPDHAyOgWPRsjie0Hc2fCAWFKmL0xAblX+0Kf2Qe7uGBMsI/xKhWPlQy2sESudTH0Rkksy/o
3Oq7M7WTMXIJ13ZVK25DHxIfQDVNtbRzpoqTbNXb+XNo4AofZ0G5ww4YtX2D6BDQByGkSNhZHmAc
iH63kd7fkvQEdNeERYbTQYPx6vNwVUWJTBrciVEzRYiWf98Mhss1i3ZOoQsL50nlkM/iUBVlky+S
hTDHqfY6REpdJV+wglOW2Dsb7FbCSK/haE8zdgY4TsYrNiJtkJqoL0IP4GSj1q9o2e9lmhHeFjyf
cz9Un5TZbPSzVAWZE4Qw5fN/Fv4T1B8iOEZXVEritQy9+xtSPRU3U56MXCOuGB+AGkgjx3j/uDzh
nFlcwUCSktlwADBr9bYdNECKFhwQ2FbmJ7ZO2az6mNhKee3XzkjDjoy1BD1nJxfWwgrm34247goW
hYGWmp4Oj9+e2XZtc9bq0i3q7VEFRjExcWQp0TPDV+95wiMTH9HgYMjdYTQ65D3gSEg/2I+p7I3s
ueTiMFyDyN62IdGS4t0BnVEprE1f21CzvAL6JQfbikQOKm9/WnhuX6viHSp/L4VVG254B4qLoMjG
zMeyUlQX7ieXxJq+eqrB45SnztGMJDaD3DqyA7hjdiloOmnSLMK+KW2V1yhiWwxPU3FB5ETW97Ox
O4CohUezUyzmcSCs1QgfaaXYywKpMm2zyEiwowrdamPPt7CVT9inqTkanvRO00FBAJ4/IX4VcqKy
PgtvwZW1V7u5wX/50Ul+IqiKeoNhedaUBbR/gsjp0gOHG6iQP6Qybb9G/DNniHGCeCXCzk2qtN8x
u41j38kZBCEPgRbEbSJNg8t30xbSnAmcT20gsC8L9UgENwzOgmZQGgoO9pn7deibEGXMPYgNh/Dr
4avBbEnPITKg2RRFgnhe8HA+L6gRa/Y5bPM2Y6W5u++nVuGrcqLHBHLUyrgXtysFHPxHsnJ9JdvT
QDtzSJmthZhq22ld1xcVMv9/JtApCAB4QDoeM1WAwEWtJX7WDhaQKSmhAA2KiFCwujxhi92wroYR
Ji3H34rZbsCEPu1gyJaBexlmOUDGVxOa2E5VUjvLv6W91tl7wlNYPFpuMsxBgow2aEm/bEYBRM6D
LDwK8ugWhhxZDzK44XvuA3IGDU6EHu1k3d7W23nBzcqT6JKnxthBgACAfWdHJsOYAJPtMF/mLA2i
sh8gR0fKeEQbOqbGEsXR1O1bebDbA9Je24H41EB/HKEtJ4hi0tec5qIwos1AmNqEJ5QUuQ6XHVkG
0E4iycZ6KZF/WF32ICWy7yalwk76ZyRcqT9FBbktChDnRYRbpqOJj6byxSVVbvD3fK8YWBYM71wY
44HSz73PenI0kkT2uD3pAWYNFJTF6KQeMrblyrRW3MTAaG9AQD3gc24J7+XdxRBL7SENs8idkF5K
QwxopBapZt9o4Z0k/i6kEWlybfoU9XEndTkzP6D6csVj3dyjupEGYsoQ1chObNwcy1zJoi7mwL0U
xwtGPO0+P1Qn5eUV02BPT9TKCHI/SAu/HhdQh2+lZevyDr/lRLSQu7p3ynViD/RN9si6uOzYOtI1
GA4ClN5nAvknsSEV71whblttst1GLSU1qKuesBPr/Cersy92IVd6IGvi9vvnEftQrMEQEHElPjcu
+YOTSzVneUjGGUsCWOcsEX2KNUQpf329kF3kf5x3bZnljKsAFV5i2qRybpR6F/V7zJzio14c1S32
H6DYV8EoNCSdzkRafr67U4bzO7KaxIv7rBDjD0NbgV+3o8rqB7WnhVylKbP/yR9YIS8kfV5HOVPK
p8y0Funo2ShWprXnXjzKB1X67JFkW2T051mtGxZ/8trqmOyL0d8mpVip6IGD/ebfSIm2K8a4YXh4
zlhqA1OdaEuweHEsgIYLyEFCRRUUoGPtOhfDvrys8V3+MyMo9aWsnXVhqEa8S/DV33U9O84oF3Cs
JtRDKx+0TNVnMuNLxY3q7FWO1Vx9BeThYkJm3HqfLSKhAxEN3xaYmzO4WL8hMCjGvOC2EhgmB4jJ
CliwA3jApzrHD6WE/M4fwnDg7IznSqKGZ0eYyEyGhMOc7ehvbeaq9harDGWJBpc3Vf4cCUFKjwqn
CctgleZi2muYIQfTKRk7J1Fhxb2DoKfK5nK+4MoyUDyhWgqTlhKfVC9wCXIxyYQ5czsjAGv957pW
TtHedDs2zU/q8tstWyeJCwCMpmmiupqUlj3tzwIheJ2AximDYjFaxrkt7usaB7MKrIvdH0cKMcWu
zFdlmzoC+kJtdqIZA4kXEW1943xwpDGB0RW1MKyhuZFgRSldfZ2chk1fBuoV1whgwNL6vBxhBUEw
6vNHmao265uCC1lp0n8S0nAg5p7W0Mely/y2x+QrvPJyMl9eIieZQqi3uJf+kHWOx0m4EvpaG3PW
fTDC7EJIZ5KYxrs+Uo3BLF3H0doGVSVqJ8upda0ZM/OXFppkY4IWyNakY3lMz9Noh3LqjGDPfOFi
g0vetJHZrobsU8TVF1rRF31AMP7Oiin+myy5KWKPOSQ1F01KAAlsso+I+TG8YASliPNuXa03+kDC
/0iL7P/Ru+/lm5E+mKhayLRXBCkA63z7dM5dxuJcodWpYdluA6aWwSUm+xqzNqcMfEWbsWWfcWRS
l4jn8eH/xX1IEvm86/bYmnv8tRCb1HTlErcxjBDM9/u3tVh5CunHqjup/q84pu/YM7mE0J0x8D8Y
8R3FRggK1wr8HyDpFS5hFxYo3EjSqrabzep1hbmaqSBmSF4L65mMxAUy5Mrx1S9PPni9cXb+c09R
gm/4lEJ4SsAeN/pvEddKEs5hq64lzbZdSkG14qj4dkBu70deW/JjtruZ7AHLAG5NFWLvfj38kyjP
EDOPf/awyIrJrpBr/LUeIKx582kpkwuexNZo54jWUzwNVHcUDS70fWOudYPagSRuT6zd//n4YPQ7
vy1CoiZKrxZpuXRbuKEBcoPuhA5C4CuMqTgnbPpJUYi/gKjzv4gF209HCn1+0muIIPpBeaIWsfhE
oToZDMA5rosA8sgYt1TQCajlbiNeO9DAcj+2r5sRUPRNYlK/XgLeUJkqkUMhLDHoFTIsQoVAd1wa
0R4lk4AWkhs17yPu0m6UnmXGZL5g4Q28MFguOJ8lyM2eoCmFm62Zs8ukJRwNVoeGKe7aiEGl57MH
mJc+Jfqc31hGuUvHDBLyNG3jBhV4NILV7hiYZU7+f3CqQ3vCz5cCXn1RPktHnjcgDAyp9bf1ugGN
NtvCnojYgN468LHUr8dULKgkFD8JiGL0vCM1+4VyX9nct29HB/dJsJ5PsyECokVo6XbkTM61+md2
o6Z1rZEItxqlS/PY7rgTaSjJd1EHOgQodays90AdCEjUHaNCSfq178U6Z6BVieogSMsTw78ruxeC
JCQ7mWLrYGIfVEwPiyJZ76l3J/wlSHy5ZWysmBlxTgyOLX4YPXJwv8cIrHR4COfn9wRjcP+IXNkH
KpwGPcWalalkacQDAQroVzOvcMHFwoCAVaJ34ZvWPq73BJ4f4Oi7J9G/i742GwLfnFzmqh6qswjs
Dg9xa8hgYbtMmq0qYP/iOxBKJldqG0X3JOCPv44kTG2lim8/nKc3/T5COWFPUBPUX76ND/34bGn8
WiXVT3YkQ3os+oEGKGXbCvBF+g+YEnUhUrZYSlbly0t1B6lzWCqwJ2mPcHrtna8zlyCRGVVecK6f
ZIBFZ9c7ycKNYTZedQzJKd+48TMe3V4D0aW/N97TKHqjO5q1z7e7Qd/zX31f7sPGAEMooC2lCQmx
V/6LZ2gt49x1tup+9AuPvswvxE7amnX3NSb//WKmY+kgFcfn5rxOBaXEgqjpmSsAUzk3GwAxtJVf
L90NjDUs7hmeZyHxD1lSYBH3kP+6fp9TFPdTNDk+/k9XLl3k+ZD+NCNd3cQR1NqtWBUTtMYez4lH
VvJ78iltPXEoc9S2I1C+e2DRIKrbKo3ktq4X5wvfvg6cI4i4zJHqNOuCoxMGRmlL3JzDRcI1kIID
mn9fZZvB1tY59Chh8jhTxuAqqc03Ai+lUAdYRgoUdY1Wafku/MN4d7DIqgE0l90udadsW90n/JG9
eiSBhqxHTTpOZIvGxxKiWR5Zd9gnbC3ZpTVLL07EPp92dL9IAXoN+/II28FLSqwdn81tesjZdDTI
8GL2VkIHMkaUrO5u36vE07NxSEYPzQM5cyO6J4/E07sJk+CaCxIRZdxi+WFgxU9fMVq30kLe7+4o
5xd8uTxs9i+mt/xesRcluWiFDtsklaeRtO95+R9fDWC3LVeReVoE/goSVgiZUTsm2xFtvKMim7d7
PkvL6zx4H9O2C0g5x2YyQBfHL47SDN/6ROG+Vq1+Z/VrDf9uHs7dmDa99AG8Kx6n9cf8LYex16tb
EFoYvHpAcXwPYWDQypFoDa3uSrdr6hmRcBI9DDo796zB+3v8y5rZtuM/iI9ObEToYJ6rWYBbulzg
/cu47KoGfIxaKCes0mLv/wynY7EDIKLYL0Fg9YTubLL15cttxFMqfb0yHBJz5Y4G4H3Xc7uAQVU2
aX6iPgUoWPO18Umb6mjqzAwQi/IYAxRg9QET/ymtcAvrPMMnmovyYOlOUx93tY9QfVyYjhXmMC9a
Rkj0GEEszXb9YRDG4sHtg6vby7oo4/zXCMK9fv6RdwJQtn2p9c8Ii1ZDpfqNhwmVfzKo0PRzPocY
SP3fr7x0692BQIFW+EB8orsog5RdcHBkF0bRGVN6sDJD6Nf5JtLnFYmv27Ms1yqoHkhsF2p6pNgT
f40Ryq/HqyNyLZnyk+IPETamikLXhYP6q4lmxj0K2hYgUS6/B75RHmkbps2ySbEWCq8MGFW27d80
z4hQG7nveKQVtxh/26sZObiRGeIq7Te+5odeAks/uO5tlKpO8LukHOPnZ6XOE0hP8w6D05Pcma5D
yFAgjG/6zPo9lRc9OOG7wuNGAcfEWMA/qP2U4YTH+t7zZKsyN3maTF08icMYOwNohggRAsX1Rh0b
hQ7jdylCjqoayc3zeorJalV48wAvcZMTabsMBcTvHE0sxM4t+ag0G2AFu/oHfIJILaWrMj9LZu4+
pnZJJjMKibn+j3KyX40O7Mc/LhLpevI5pyEd8Y2fh7STKUTdLY3LxpgCQ+6g9V4AaVFjnt0asy7r
neEUdWNT+7zwFtysPpCpeqqodiAwENMQ7PP6+fOR7iRr7QwzvJXiQH/Vi6luEfc8+EeI2KITtO+7
1poMjdn6ivE6T77156N/wq6dS9u5FGgX0uljtxNZMJSTiJRXqNNMd8s/LAoi+xa81Wt8+4kamF3p
RwNFnnncGJCvD+HWXhh7PdqsRJS5CfHjZMEKyVGZ6y20nZC+YC5YTI+rYqtfNrH+AIJhBLUTIufI
PTfcn2qU3tBkwjvuGmrujFYA7sbC2NWGKwc8GSUPMwVChoATtV1DQutezxbre03+5RV+ZVZujowe
1N3TxhKExfRzgLR8VuO67Qkbm1Exl3pTl/nxyK3d8HGvkhHnVk2/LMfo/EQSdgUw7V3bfGblYOoW
64v5TyFRWYFwGlJVJrDeagn3ZPgFCqLMs/a6u/xrr5uaYjK1MR4dpCpsudg/7WOCiRKBQm+xapIL
HfbQm7CZkSHDaRGkY5v3befvkVchuTQSVOYtiuJp0ViRSCGbbTktCuKRhfZdK9shvTYXYCVF1JvG
EB6+5TJUnycUTTTlmO5WQ1qajDe8vx9WlahbwdiJiN7NNw0I5gmLgTZcqmyDSqeYi9HkkRvy9JWa
zBJAU3iE6YWtmt13eTvjaJSXGo1i/jrQH0yPZNVZNVgUltl0wGvcNXXpkxtPCEXkaSVAjkRUo04t
rh3L6qOt6PK90np+lnNxW3JS3gpYvlIKdw6nXpvAxhhfbsncZLMaZSK6frr3Oit69vadXBRPW7Ih
1Vnj9MUiCuyKrJh3RDB6Nvb1B2aXsdSEn3Kx76oBGmxpDmvvopSSX/LX2RP84XIW2PQOf7vJbpLa
RLBY7pCAhNSHcN8pzsnSMouQAopxFOkEpiXZqPZ3MuutGkC6wmDoSwn/Zq2OBwK9VaZQohYfuY+m
uzw0IMXhxuchtXo+YbEd1Q+dLMdZIzY+ZbTkM+K5IkUFl9wOP0X0OcWaIkhLZExsNa0ieU8O90Ax
9TWyZ/Wrkt1gyl3lxylGjrTJ7YzlEss1H0R5zVxY4cEsr+H+u+zXeQZQw0v8zJ6iVHybdBb5iBrA
DW29TFCRRbZK5IOw4HlZIxBoE1hoK3iK3OjpOEJS5X9ZkmtYeyCGdpkRTLZsQN0m2PykHo//DUs0
HIN+NcCA4jejI0tr5KQahnJL5VxrHAiqfP0zUqlJkG4XB7EpmVCo3Y6iNGCR2NRJVmoxNBSdK+C8
wiNHBWSuzCw4drkA6Qm9GM7lSh94tGdhKXUsuLXc5qGxYD2ZIh5Nui3hazmyqqwDvKtzcfDtr7u/
P2kqCRuZYQ2NLF9zdFW2xYm4rSXh0NIrOEtYvi+kUCyvunommOe1gPHMbq8D7Qv1vLpD1Z/8BrNa
k/WdgxeRlyv5fkcEpsKJhTnI/kDRPmI1MJsec+Q5C/8WLtCkkbXbScTB8DZiiJ6BkosCiWjMB/QR
AMiGfUeVIXJYvIzR+26n2g0BX0zmBGhYcux76asOABZFibK/ja3NWYIN4saO4y3QoarPZX9VVkXy
9j5aNsdB8KxObd8E6LXE0W7fZdLgW8OhwXKvPX5YoK0r+ITpkyCbVgJlSKZlNP8DZIlHCpCb5cok
SmcJWeD8XT5P8ZgX6cDgf7P5FwFH9G/DGtfp6yc5/4ZhAPFc+StbTNZN0MQCwJh7JSSLsIogBOxr
dg1Iib6CWKDrnPE0EXxy16Y2Fjht4zMwE+nGW/Ssyw/DB3+rrra3C2sz71Vn4MYHvgsmrPQESF9i
mseLvhwF+RqoRZanqH9rI5o794+A96cglNmPZ3btS7LZaUDN2mppUeAso7MTSzurQ9D6gRLtXFEZ
/1JumSdutLIVJDXLGk2IUtzywsZmltYJUJubrCp2xbT6cniwRfuiNC5A/aTEDy8/no1X+LN+1IHc
UHVPzczjJ+K+1rvRi1ST10KCkThKRvbFVPZjujigx50p52tXQETpEFQbM+fr/ccoYkHH3e7hbEDX
R8Ig5Y6h9vWwVO49bBX/9HjOl1RhuRfRPlrQvBrMz3babL+09Bo2uYDf9daeureYdKYHLqfIBMjM
tHrdpnQnFNwEEQa0NSHzfyQmgRE9q2SzqmLPjUZjYVhZJC9ofzNKnN8E3AtJp6jsPvEByBGU9Hfc
mMFlfvUdjsS916ubrEGYLxpappcpny04DtLA08NZLz8mBquaTmtloEGr03IY9PAWlo3hqO8k8mle
xCx2W1o3Eun2QsCQNQd1A2YQ4A2FzRKYLCnN8BJrMHw3swLeqJOiQm+yQ2OzAi/PrXe2uUpbWycw
3+JaCnaeYihxgGfCA+ungxMRR/4n1XiMYyPtrabte8fKn0eWDi5BjkgWy9N7AnEf7Vusd0t13Nx8
LRuiTZBpfNK0Af362CLcEkMZpY39q4m/MXKZsvJXPSsUTeo6Yx1XFK+RNanB2MQIwWKs+i6IYzR6
P09XOb9BP7YGN2xDk3gGyq9DRCjCD2NlUfsnzPktgB7+sJTFaUESg5OGlIyHpbO8BrmGGVAB0MPY
YJsEKbp52non0UJ/EvwwZ6eWpQMquOYw8IKnqq1LFuNME6F9qGImzzm5rl5WwrbsmhVMVHZTsD30
P4TGm/hmnDumZmcxFqkhnfHB/fN5j8OopTdCHq65oUwfUqI7RwOiINK7IfIhbottxNvafdTmCmdG
Mb8NjKwvo57ynzD6EhpT3P7uaMUWWdNLtEDiR6aqfLeyQoJdQmCgJX03AWqDI8ME4Lq+KdGwoHJS
CcukM0dfiarIpClQtZl1PorH9rI+Rmeu7VzKg33eZFxsxLAcKqmrqYfyp+jmS72M8apMy3RbYflp
BWU11SIHHrhKeLMDSQsuL1tnv5rUxBORquJPLkj+BHmX1sQdUkyyZIa4B9bZGNEKnbVzHLVYEztB
GEtnXgUb3UVtyQDDo9pqg8HZ97ipJ9Oeq8T09xP1Ekd1WZQxda17Kt/EjFHO0v4xGTa/AR7+xlST
un8R6rFLpoDR8InjNHk+jJYZu7Z78Dil/wxm64Nt5MYNmYbJE0UMADomSxL9P0Z6eCMxAXd929DA
2yMsfhIEDVSqfQw163qE9d0DVYstVd6WgFf/l1Fk2HEDR23XEps03zK6nDAlyFEEAGGI0fygIfQT
HCDcq4fG6xb/SF1w9cUbYnsSsnKATOTa3sYsKCW9DmsfuXMBLybzMfUVuy7V5Ac+FvyGSugdLah5
19DOqyCIJUsLhKwzqbNIToNpw8b/RIupWLPIPkaLUCTReVxyGaVSE2CejFtiYMhUBUHDKYKZtwKW
63lIVC2Tvh9P5DpZ1F7QhRhKFO+kw3oXl40stksKxdbopaReG2IqwWamG30gO7bJ2mVpci5n/9Y4
RvRJGwUavmDgGvJj/hGFWh79gvy/464UNdY3Q67jJHLCuSTfc5kwrDAPJmMe/IszwPSB3B9Sh8pV
sn0iadL+31W9yel6Y7zIUwn9GN5cnTRIZCsez7IR/wYRTDefB5LY/OyGO+zscy/tV0cixVLnnUwq
veTAyxCuJB1zHTfetjfXJ5Gi4nNTo33+Bml8JAfrwYiQlR0ICzsQf15rVwr7r5pI/hYeSNOi0W8y
HeXM8oL0OcAgnfcVeiWgPOu8qQwEKlkjy48xd0Bdoxue7qa50Irl6JircMPwZ0D6ZGfiI4dGqDeX
RUM/fcEDX/pFGX3I3eXv2uprN4iy+Z/24YOMj/fFNYNCkTdSvgcyguXyr9L70YfXMxxOGb2qRJuN
l0uaAocwVYngGZhzZN8w/uPNKBCfCd3wvferrimlCU1GfeELi+odx5Cc7xtz85+ZtVh0QFZXta+0
W9DphE4CO1eZSw+JB3cREAVfjF33JXPknHO+Z9sib7ksE3NoGgd5pAyYO9c498OLbvqAMHtwaGws
a5kefV3tCWen9bYQG9P7cNHwSHGCVb7Cbflcluy3J6HSnJGDoid0jwI1fZr71vCPqLtZ0Z8aRtXr
4wPXc6iACmq5cLOcIC75qNFOSrrq+hFh5u8Lv5+AnCWq5ASV9vDEYb4tL0brn0lWazi1JvWPERq3
8q1hLdfuokSa+1v39u1lRSiMNpeY/zb3mmgU4+Nbl677PpUjNGDdVl4uXrXvpYBDkU7SrKX9r6fU
nynM5XuCybS2AV+NyanHNH+e1bSyEWeNOEG6enhzC/Ap2Ff1vxyxBdAvI8/9vo/rI/r0wLy9db6t
iNHwOgVIUJ/4I+4a65uRe6zeAF6CRqllRq1RS76c5UO/jdnY1Eg6HPFZIhKkSWXIgN3kngUcEpoU
VwmTMpmm2jC8ie67+/+t8+3xnnDzNJIwKe+M2f1ephm9v0eELq+kjwFf5YY0OdOoEZrkDUfIceMF
sKwthlUtaX9uj6aioM5z/ApmwjLHeIQxL8JtMNWrU7cttaJVjmkzZLrUf7t0kJIPXLusA3poAJrT
eQTnDCXA2LwHZzSAKEfA3D5UIGuLgpbRMUfTACxJeGEIbSD0OZ18zC/yWWMiOaJydYq/t6wosPAB
Rv0jpNaMUUm6KS1Gg93gv397N7xw8U2kvkpbeIa0dBXEQghAH0Kj/upihBqu3ls9OVKNC1bLVgSA
G/UaK5qJIwUzlT/O1Tdwp2XnImE0+w5ZABYsKje+Q4GddNAx+33y0f4kljnU3bILkEx1yoTddryr
pMYggmvxpnPO9KsqoumOnPHT3rGFJy5o/NtU/ETlIgrDm4+ZaOj4qsvLq+UGYjp2k0M7XXu14vfJ
OnIlBdUHOBDG9p26bhWgibQC/Wp5gSNGbHfIRuAE5iZZQ9chZhZAkVoZ0zIMbDJXR9X8/6x5e9Jo
DtPs5P9KBquVXQB2tHNKIQlBAMVxowoU7knW5lVnsxIC8izCTp//sEzmZRcszoyw3vyLTycZsp+N
TN9Ep8c76X1n5jVXmgXMNpvr6m2Y8Kq72zHtpqoq4LIkDTWx+Sh2aDEg4OL6AAbLuUJLsm5NTW5u
tCQyPpunSZedHprKhY6gCFzcIofM4sR3/lJwa1iRssZ5/CRA3EDXYECObnBINoY3N+KKoRE0NcbV
aH6OI3JuQMXJEz7Uyk2Lu7/rwbDyoZqh1i6ieLXHEZjKAgzUWxyvs8jENFrUe9x/MhxcnHujShrn
vd0ctq9iG04ixrSAD1EzeV2LZG7nYJcXqGpR65Uz+wYrNw8fDIDaV/35nTZRNUF/m0ie2msvhocq
akcnu1QcHRow1Ygu4M/pvwt4p8g3LmNATep89A/0z5aW7VYjL2+dHDzgSXQLzephNyTjyLIAUry2
zX2W4ktJJwKRCuIVnKD0UHUd2TxYnEFPxEQPiRKQNVcS3ES7Wpj67CguWQ1r/qvHpgC4XOADUBMK
+wOrlXKM2WHCJ15lqd3ghLmCCfoxy04KHQk5LdVFT0d2avjz7sAUaipbxJ7Oz9cnbPnhRcD7lei1
nUTSmXolpAcldXVJ0gl/NuZM5cUZ5GAtsE4oRLmElS6qZYiuP8zLPRCvOXMJGxLuUMMQuPC/0hVQ
4hbeDhMD616ehpjmYR5jgERX2zAE64Y7kgPTZ1nUg54OKMNUMcFK3Qh95WmwLooDZ+G2cuKf3mrB
82O7Mbe/vYelpr3dKH0onKAjUMfn2UgU8ovsmv8lzgZHWvyqPadjI/VdjhlJtQDg9AZ3tmjFG5Kr
r+aTSSQ1og9qjRFIJw6eaksQ2xjHxhjactCTcydscNM+SGvuQ2UXT1WvN1hz3/xHK+Zl85T9wAfG
GuebFEjFv0/dQmz9Nvfz6zgR4qhBJe6Y9oPH2tb/SflZKfwPvAszJ3L7fmcw8xkfA0VKvwCfw3dT
bZoX7rWYw4e8nf7fi1vqXaapDV3u6dRWjw9lsRBwXQdqDKcju0Z7PA/FG++anaE5z4d6ggF9l9GX
mKSOr0f7abcbemr2JVT2FnP3pvPKn6tI1Uf1mmvXRxTE+F5mMgO6E8Bo+T2RxEmJUl8oFY5cWMHZ
+53lQ1vdaE3tW5I57x2qySPmtXQ+wFMWumddOxwH7REa8yq5sYnd8Ziu2gvO858Umotu7CQwvjlp
XR92SVIHaMqvVN/38opkN8IZ+LLbsj6Oei4FyWeP07SLsiZCX0N70AeMff1xz9954CfnAVu0J+3p
NuVHyA6uWlKIljIbthN2NKRL8YnKbYeTophDIv6tpVzoSO63DDuWAlglUUL6WmoWc9moVFJhSlGZ
k8y5CMKD7t4JcroQwQFpccSMS1PhhIdsLzT/qgzK0dEEdZhqvptNQY4H+RF/f/Iyn8DBEDqfycdR
9Mr2d+4syjWzaL9ibBzKbacQegG2BKPo42TYhmhXYv4CbTcJ1IXDct03s4dxgdIW65b0RLZBwuR6
9A0rUZoj6vHcUzFwOvqMwaLQAviu7voSJJR6+SFr3gUu51/fCziX9MogxoN5YpjiyjcUynv63y+u
sD9Q9R+g8jrKQtSZVOESfh1Luhv86Biccuo2/Ofs5s4BLO+zPEfV3qrvQbJyGU2h3wxQZAU9R5yp
bnGlUE6cm9Rgod0hQRCjAnCrV9Nt07bmdqOGZFrSFnjYrsmeBRYZ+mF8mXF+Tf0ImU8J8rZbWRU5
40rqrBkYJCMB/u78x5IyE9x/cKRjtBB7mYYNZkqkXA8nLSCg4xrkYQKrfSPUn0avGeOqNtg6+NJr
0S4Xpc6Y8Izeszke8pw0sGsz1xZMO/P7zm1IwM9v9r+rg1nmOXZM1HqMKOGQXHu11K0pkL/Hpx94
ZIquxYOaZ2EE5iAZWeAy3S69VW65mTveqZBfe8jCYsYL6NHmhoWMf+406GPD0IqIwxv1me3Z+veK
zw3jLKHn78CzPJ3e8W5X6CireSWBrdLkIi0BH/AudT/0uGi3JSs/ZV8M7HRyWJrDY78ym6+5twey
A0FqBV59jYYpew8fpHJH9gx9Y0P7jM01MmWDkrMwkL/WYCPEt3R25MDktJdP6Hnei1bdZSr1vnmr
6Qc24KTIOguC4iP7iz9EVbnDiymOgLXAuoKxRTFoPWJddKXP2wVkyX6YU0YsuxeWfc87gg0Kor2m
az8MiaVlxLRhewRVX7pIRXEIIaM0MVQlMkC7Ub6Wpt54lNAqJI//n45Q7EGiryVq81CvMx6Dnjz0
yrRqJYN1+7MtaAYXOwLQphvXvfVHAaAFLveDdF2IQFaux2QmojQEqi5e8+agQAnUE80AYEfCiy1l
7nEGmLYQvyOV8c1rPWrCnCvjE9Mwa2vx1CsfctL9mXtDdHGuLCSAy146eLg9/+g3/UDd1v5EePX2
rrAaRZixsInLSic8RE7AcwQyyC64gUA4DKmTnzExrHT54Q/FGfA6MKJrgdVk9lHYNwkXlPxtLyLy
6d2AhONK+gZ0anE9QZpHFw/ZStvp5QHGDi8tBicbATgXtnZ9ZgB/ZNG44wKn24ySEZz+uN7NWMa/
8tnTBXnWO0QUT2IjX5Cv+jpOHa7MyUjQKQyhMMhl4MLXDRGFxLPQrKNV3dg9fH6GMYTq+I6gQVGj
KYmyeEnidDIqZXj2lZSYDIX5X5iclO1PP/DzUKAbqkqU3SxfvYj3sTGdQ0WKG/M2IPgZt05L5ExM
TI5BFs+grBfjKgpb6DDe3YRk57KHoljURe6bHsS7FXKNWrvo0Rj9XUq++oyNMf9FH4AHVNdICIax
IrZiaxSp+llFsSKfTvNiO6EukoYcBNo/Y5MxQESvNNd6Os/UD3aoMra3jKEJlT/Eu2p8wHG0glVe
fuhsGkdpGBC6BC5jgTSt8DXIGC6NLrNid78dVr56aHrMH+6trKi0g5S57u1w1J8UOteAcXcTbycx
2vpvJEK4+CvUl8exywlQecZETAMChbRyVKiATDAlKIA8VUXf61bnbZRMbMpGDe0BluinZIZhdmZL
7DOONngIo77Pblti7o505ek1Hp+90jAcNN7Cp2Jw8Zts0+CWkgajj/b2YXC/6CLJV6lt6bMqel4R
xY9cD4CTUlAFwwAurvF+WqB/ydz7xyTfVTpnZ5jRuLCpv31W0y2y22wpCmCyigEshhhO0vffKP+o
8stL6gSgoHFAAEJ1vDKu2J1iR1xdS0hYOwctUU1ICrVPey6cHZkAmW1tA0c8Y0BzFREvZ5GEZa7e
KZoKFXTUGomfkl8xIAIiy6/S/oTArHNJj0/0WjYjrvKiv8VyivWMsV0geEObv8A0cVeN3jPC/SkK
DPB7b3PgjYkzxbxAks4vS9jxaLcYvHcUcTyJ/z9WbzcZPLrmuM3q16dwpgVo/lzHZsltn8x3+fgd
8+jwDJrVVrBOBzRf9ndX/0VYfm6nZjH9Xtr0XkFl6lNp2koizF7PZw82N55SOKNgybcCYn8M38jI
SQP9s0gys/Nbk0LgERI7hu8GCuagFqHUwYi/ZUJp7JWQ7HanaRjadvIfTYNmGfAZQBNCz/ny8Ysl
x09cluobisMGJ9NqHVnyTn65af4bDxZFw2K0UP6KIEvbzAFjv+JxZSkhr8bcr6chRpmq6IiyyZqu
VVQyjD94qdYTLVOkzJbd30/abmzODs0kYNjaGNo9VRl8q/vXPplQD/phy7XwlvxOJ3xsMQZlWYKL
7vDwdfFPd6QdWTxA5BtJzAcPZIotMnWHuIMhgX2RItY1ZsU3fTX6St5ISBqVwzI3acq5qaZLO6qo
kVVABEfHy94KrqsAAxppFZ3PNetEol0IC0JC6AI2Km5wMbyvb5eiYK1RwLK7aDh+EDoGayyUCYoE
Lhkp1q65liyT/425HCZ5dOCM8I2rG92t276tbNNt9KXEICVISMGg9aV+wbjQasnaR1BPs+6kBjMQ
J5yHsisMs0ln5FhBmN29Kad0waXXELO6rKGckKJaGmG/+Ke3dadnxQtLOQQr0LQOnZs5kB/EzTW/
yhAsDeJ90u5A6hrC527Dh1Owki4PzUa8fB3QWhiEXrGsoCkodQKX+jjL94KVj5udzTw4Oiry6NSH
eGDjWfwC1hx+2kAuK/c9rvGnKw5a3Bkdrr08Ar5DvbnCdxRZqm5hPbS21GvC2l2/ikI9O3KDIe32
Irf5iGhcucYV5a1sumPucrpOdkpPAiFdvL3r01Mo5N1sLuZ0DYt2JK1grwoKUWJJa1DdM6wcbFH3
ogOZ9HrSbWv6jFlqV/pEfAXgr5Co06i+DXu2+6bxMPdanTPr2o6zVqv3Meeix4GDYePGHV/H+CCT
B9CKVvjhDddqfbOxtlcOeEQsHx1RyLi27sz/01ZGOnKp8eEAhtlffBYJuIGrAX7BDxd9jTRQOfWw
/fdEcQqjKvOHiLOcGkF2NY7WFM9h1/q6Q5lPa6DzTL8K7jSANW5/yLE9zmKgP9b3FlsX5fq3wgsp
iZM6uKcAvao43nUYXd2dgrLv1fyPhE/mut4uHzj4GPN3GQaRw5BMzYZFsFympBFD98/cWx0NGlWH
vVXM8amRSAn6cYuBdqM3nIf7NrWHf8D0MZASiLxYtPmVe76NcFux9FmKhMnIj0yBi0J2UBtrcFo5
RH6QSMelfaqVeuxYDaOvjq3Mhgp+SUBxejXy1Q42qumeoObQle6s34bCAKUyeKL1qC99z0JB+e3u
0CVqXpGiSXodCI6yEnRNPspOMMkYJM7jaPIPBo+bqfm5RG0qsu2oMZXokw2YG7yqqyzah1Lk7b01
6857u+0PXvSqn5FCrxb01im/6SGOfyzs/RjmZIW8QRtMmFdKDeNRNDxzTmZrJ4XjzS1TI/EA1z79
bM2rtbCpmyZUKyU8/PDhZ+IU8BzjAyedVfZ1GThKl2TkLlgdOToUMmYLd2dcYlEOTJU+vJ3ngTVk
L6QeqxhNxHzILVGuN760JB0rUiX9rGizLLbySwI7BMrWxvswzzlVXnZ1J8LrjnJrXKaDYdA5TIrM
/g4VC8gU5mp3tbYi2HJ7G/cMmqBz23yKMUzQSIrhg2l8Z4z3Cmt4Hh8d2Pr0EuFev1LnNgtPyywj
7fvmz2JDYV0p6gYLch08beaOSs+drzeOoHpezE1+nupfAL79F4pmBBERZ5vWHBwqWuxJywxyBzIy
Vwk7BtTEO3bdneAG2ZOqEkQoyo7jmiSewc9I8eGHkX/aPvsxFRF2emEDzR7u7GUzEZq1iya2SHn7
NGkKaLVzfDyVQhFCrexbBM4Wyui2BaINqQe9RyGNpOESh9VvuRQJLPMqH65ZOAXERHy/RH7aE5W3
xfMDcUGbz30RtePkdeWlmyuYbnAjotxvi08YeHoTqGrkoqFdr0sJiDYj23jVhAux9FEO4m2sGaYB
lU1seOzJV3vpPLiMkAbIbjC+6dCnDoMFsSY761m5t4PIvg6F51vVSZD469joBfphTrDWMNQ4HPeF
7CwcH4OTCbdh/onr1lvVyvbRp6FJ9KB74/tyQuxLwzRRAn/Il5ejPUSg7H98HJjRMKb6xeiT+veL
hf/yQD1VWQ7bgKBuVLH9e+lxI+20NV0iswnVkob7/U/HD8Ai3HtrqoJKueUtFOxOQ58wdQicRgFA
3MeDeW4PmP2xuS7lWYuNt4qwK0405tiit41rjxT7rrSXBClm+tbJzTpWYRAD68qPcv6dFOrO0k/m
/jqKg71McNnGuEb2pJaYuqfmCHWEez4KgPuhfz7Cupf5vPK/2mucXs/AbY2FNcBUOvELnaV5V0sr
qvy7pr7rDhhb1kFblPNz4HsQwuYutN4/ZMoZGt1qIOe/9PqkTtE6PTSROpCGJqVIhxqZZ9AayFGp
iDB14fGOBrDkfGOiRKSMd3gVPop947JeCquzgjo5eFI6a3qu2qFPwmO6Y+qkanklxrTLPQIs/JbG
y8/j+Px/SgIGQvLg3j7CqFpLrsFSnSerliuWYBJ7eFJjdP4bBdc+0Sx+B1peH/tY00HBpz9yHmyB
tTOfdEFZyrLgYVVBt0+NcMZvWQpw4MMb5fdPYLIj7+8TtGL0Pywk2118CYaztZZT2HZ4rPSH/aSM
79D+t9DGQWLBhPEHAFQ0BVJx5k+lKK+W+K6ur1YGqYGjaX/3XSBrUu/5Vyg3UKAKe+joMU9NMFyH
HyMJdwaAKY1nuXhOymKquVK1t5YrRoe5ISFLg/MPM0+NXRES6mtnYR+PFlkOAVQplN/pw7EFxOSr
cQhmkFLeJ1Zf5bOTeWWLXsFjEaMQ9NtE3J8Sh+PR+Dj1NLRK25L6gI7A2wpBJcouVlk41n5EyZxx
6Av6+hxGFELrc2zhz4v44hkKCwpo7vshM33JtdA1sgljHjOlEQE1XnrKwWStUInfdbJZ5kVmFrB2
Bi+6Ek7TvO29l1s6IdS9uMCxRJ6rbsN86zp2LMktmI7VGBit/S4QTuYpCU2zwatYXpRdTdVx+1Fo
BFaMQs1JAbmclbZkxsL205KnvfU0sFYOZI/Mu8AG+RxTzb3c/Y89jdlGMy3NXt8c0Bf0RON62xVg
YLGZja8vIh/nu4nMbUvBYtPHAuqnNm+gxx0RuCAJNB+unweF7+pkuJNH35giqcN30geYD+r8SyvG
RrHQ1+ihb0AWMmodACzt1ENjB2PhKtzS4lPcLhNj5/GK+qA4aJOeoARpg6Eaaa8Nim1MCKHOXL66
nkr7HEueis9QgHelAM/UNMPNG7M17Ea/KjRJVeFwbtzJAjm7g2UnOCFl/q1NxP1AF4bby9ugDtSn
HpxSosgcVj0f1mC2MXfrzUZB99CO+SL8T3myX/0Od3EsAKqvtcFe42+OmfwFVWM2aHuRQ0jxpP/W
0spLdYTiQIz04Ivd9gZL47kWS4foFfcT3LCv6hxWONnJThoCgR712rI6FnjlkFBJEbTnv6qQIjNF
Rf1aJ0Y9N2g4CXVGeJA1KJiW0y9owyJL6LFcbcuH/QHBcY0IhvoZRXHhNSXZlVLl/Ssb5FLxF8lO
pZQrun0FdSStpRxujSXuOhRyWYGmX+kfVYC2VRSbtuZG2FsnskM2I9VknNZsvyTxnayPrJJ2zzD+
BMWIMtrZOXl/FHzpPfnMVJVTg4c4n9l6slTd9jjbepcAL3o8fy4HrBMzVpJNlFsLNxXw2fLvwgxt
kYLs3Gie8RUJfTdhjrY5FEnnvNm9C0hwrhPlRCGDLEYRTK4W1uPjXASxBw84TuzI6vTdxgVs6e4y
68RPULalpwll4AreIBkquXQ6Xy82jG0ttzENWTx5MSLNuwu+FOQcnwFFUL0ymjkqV/5fPIjIX+hr
knAprqV+noWLHyjF1H0lUjxob39AxpWEl6Fgb2npl0bcLI2es+Ie6V1PBFpvz+VjsJWwyD1V7bRD
0O3ZsLWI4wRIFcWBl0+hRFx4GWf/wUtiphB4/XO+WjZeEaca3duIkNk15WSuYcEM9FPv37dPpSA4
Uxx3vQKqJTatoakZWYEM2No9Py1AUlu9eSi/iRFXnHXHk2VQyMwiw3kslwxQBSn/dv7jl9WpKyfj
FBCuq8+5MS1puPIS2qoAGNctLzyJUirv7FeSWHdP3SVvwjfeI7nX5nvNC2G5TB+sXCXIsC+LQbvX
g6Zq6l2LwYTGFwfOmSxWF0slv/vInHVcU5Vxq6/fCzYdKCTiUYrPBUa+9rOdrfIKbckdL73ox+sE
DdtD64P6pX6crGNy8VHKuJ/qkkBMwRFQGHqsB3aX/mjUm1bHP19CHpTDv9nLm8XXVYiLQHPhC1IY
VmCK4WSxvZpgtsF+O6cJ5kMkXBbD8BQUYOJJne0P5iVg4eKowcpp7avp83G4zjlwWFVP/b5D8w6a
MXlpTgBcZk95ZPGovPchaDOUG4S0mF7PvclfXV6Eqz2eO2CdyHQCyKvgxEMM1XCoewRBARohpFCR
lfMdBTHQcF6UoduUCG+CzucgUu8ZhLPJ+I5pMNro7uwdtsg9K3datlW6+KFwpeN9Iv8WjWB9I5QM
s80WGqv82OtmbwWD9Gv2eVSCErDry9cNabv7818g2IRpgtc54KEl5GDDTNOyBbltksRYogBck+j/
2jkl9c7ZdJsqTtuQLQBBzaRoWBUb9rcKOC63SAOBXC9jn67bPyfUJPtd+Xj+UlgT1LIohYhiwxrx
0pmb6685YpyGPqc0nzw6bgSWduTlKb88GOeNH5AqGVZI6Nb0zYjH19PMm4/bCW6t9kMJKqbvz8va
eOplPQAfI6aGsz4OZEaIM7h+g3/yzwOQ8iA8OLR9Lss44MrqOF1QJrEpewfbPSKL0dwVBmdMbBFQ
zD4uH8pqypyiUVY3qPdao2flDpzany89YVmYpaspMhv7JOaZhDh73zMwELXTSikgR2vIKSWemCRC
Y7OjhoKAwFR1+/kqqeduWRshkVee9H/Nwdn5tpkD/yK3WKGDValfdRlnDHJyoEcxlKER8wOTQfgJ
jo5PUU7tHd8yRAu339sh+X/JVIev63bSZrPLcKRhI/xQYGZJZru3U5Vni+j7pWNfco4Kq40fd7ps
Fdd+eCCzPxm8gQLtoaveXwVf5JMokOzwqi2AZZKQSjlbZ199dXY56OVKHKghhPfIN7iSQXSdPw2u
feOP5b7wPyHRaPerjtZfGPyu52Hdovyx12bNSMsE+Fy6yWfeVJKDqEL/b05BgvLSqHn1ypXuA+/n
CfsMjGBz20C4Wbg732Bt63aM7fnsawSs8L17hq2kmxkHvmsCEP8buWscg6sTXWVkmTnr11Y6LfZy
cV7RiNvb2+LKiiezMFOXa1cRcDnwOqCGsboXcjYOqZQY+7gmlbalHSUQsdNRsd8AXnDVmG7TlCRX
LAhKCGTwSHxGPOFZnB7aWTPVh7O8MxIvUhC0dkIza/3Gb1jQyFYSVDL9JAMO2bXEQspOPXB+dgUq
XT+oOOIpWsMdyW8Ixw9mv6xObfYZ08Ib8COYEB1ewZD8XYRsXUJOQmvpdEgEIB1pvG6e0kkakNSp
MPBJTYi1KMzCYWvA2A3Wrjcpu61zbdzfY7wf1uHJU22ifZm/+CrHsGI5PPuBqXNawxgn4suQU6Wb
g99T3dN0qYL0rh8ACLDz3mrkBY1LvU6mkiJ9cXNUYHQSNJGy6atHb9iSBAcUQr00SPSAU6GVWSIM
Ap7n36X+ORv7f9axha+Mgffcp3glIuCOKDr/WCCP+9qaaHhv+bPx7C/r9/pawXKj/3vSetGLX6EL
axcyCZGYYF6JqSzk+Z5XMqoEGztj48ELGywn8X7LzRTNGum2jcA7D7zRkn/QiGm/Bg20Wg1uT5qj
QUWeD97IvEux76N1acfBW1eY1IFtcQCW2RKzwljX1VjXVdIgm58XCyvChQzIP+H8xbUWTsxJxFya
FouNaQpZvfrC3pPflpLtgJqZaezlvLsQ3K54AqN8LC8V0ysOr6AIsPexW48Hn/9cCYxDrfRKmMRX
yu6iaoT79F0hw4U9Mac7+F4IRp1f3b0J1vbMoOiQn3Go0npsPOtsy6FFFZXyyCX+FPwD3M0rmiSW
zPnlLw+rL5OTOT1ofviTa1Ovfl40UB4N5qch1B6IimvzrnnNva81XaBN8QKXdlJdFMupz+VOB4uv
k21zmoZEGn4YIPTQHLDzGZOtY5ZK368hCwFrqZDvIDqpnrQzCbRicY8ZR/qdsjMlAsCxk1xeSnfE
Us5pxOXDj6kVT7AVf8AicgTr5FvXxzGEPPeGpC6yxpn0zGHXC4pYmLcn4dkogJy85gUT30EfJn3V
pkIMLJjaLFxDcnyMwZlXnfgJjSMWC6C9/9Ik+EgmB5HYo6lwLSOD451uLsJkJ+vsWy0G6kUK26Wu
q4EpEACREz7KqCS0Gy7MzckpCxJfSXQNFuEM5hw7Ymwn13upq+LtNkLkwaG/uyB4W2Y4fQo+et3y
gZtdqud0UHS/zwaBSgnRWwcMrgrjM/i8rYVRQvBaBHdVAdT9Am32WU85WuAqtpR3rqSZO1bZP/iJ
RqNE4LGX8BtOc3ggH6EddUHepq4/luyjQixgNHVjmaG5EcpuKJG57gf8GLbpMGJ/RM0FtMjIRRrC
vZ1hHHF32pRabPoNwXJZnwzangyVw8WTfO6CH2IKNv0ctnW63T3y/AZKvaNpLt8jhzqiqqfZh5Ac
fgqdXWEjf29m3Vj5sP9j5J5zMWiDWod/y3YmMbSeL6eKioA7P9j459rQQEzBI3NzsNJ8Ki2pY6mQ
d4gypjOlXsM+hWAzoTNBNm5Ej8tTWK2LnXRfPhO/X/uAR2NuIi0xqB3Rk8lUFfh9a65hp5nSnlkP
wUsCL01xhN86y09mBsZVgSkkSuwjRFSJWFmkizbba+xvRTYF7BLV+pCcXhruhieRNC7j9iCouHx5
JNzyL/2Kbg+1leYgTKQFjciUQ7Yhbj1tzNpBxPHrtRa3O9OQLXdq+dXiOCPy0TjGtUMb4qTd926+
WcLYRVs3kqUHs4CqtdWVEKHn2unc26LulgJTEr1H25qJC26fECsLeLRQld/9eciApZM6/3VNj8T0
FbPKRnNNkaAHS6V9TUGIi22BeZ23OwT/feUIMwcwngV9Y7e0XgPQxQzG8Ai8Q1V0ss4ETphvmeqR
mm0anyTD0k9a1eh7MJ/916k8kPh+k7Vv0ukZsCBLzVrJBc/mnEJj8mFWqPlT8M/e11v72vOKhpIh
jT9WOQTMywjUdeEcV1aazYbsFyU6DSYjewd495KQMnGHy8M/MVuNjhRjfG71DrK4akd7fqoXYoXz
CuiNeCYjo7DeJ/yy8rgVlt0/X55Zt3fIf8MossycoU01c2NMu5YHFL+5x4PBRS6GlDbWNcP+DFTL
YRVPY7Y9/iCZNH9/4E/TpAUonuYE7xTSOdOKK/pdFePfuofJiZYs2+i0RpQntPEK2R/7vpMTg3O8
iCxFj1ABgLgREJ4yg2TIPXVAZ4Gm58Ms5ULaVNhGF9n/KFuXYdgn2YNJAs43EcyiniLn1kef5WSk
bZawPWIfAp4aHBx4/cXY+MhJn+76WcM4gtXZhi/vNcwzHcFuuBVH3WbhB1sAyYFdQvFMG5DJWsqg
4k17A7nuRQt9XwLUGrKGVyyBPK77U5R+ChBcaZhnnn970s99QqBQdcLUFCbA3ElclHJXiG+l7HTm
cArDLi7ZArxKlr35+ZZCo2GLsWzQDi/91gjCrg0ZV2pVbB0XuSLGmj8G+VhI935vJjyuq5q/lDxK
JMNrwZyfRML07x2jrC5xzZVq82hxfGQE95QQDMrYi4r5xr4qVSinhuTDAKNDj2YXFaKvj1Egu81d
sHb21llcLCyLd/1BSPkHPPbcqRikRvlfNTVCbK8aar13ArKNiefUAqRsWI6HYeRD7ZO9hBC5kfWo
PfUS9MCjI0gMlY6MtMcwhezhCa/K7corbq+c92D25WIPWKta7Tm21Nf9rp77kgO/qeLf/57isKls
w83EAvHno9YevJkjoESj1cMZ10VAAlWJtGjVLQEa94wvZzn9ZMZeLSzUHPOnpIJVGWGG/QLIuiWt
X7Xuf5tQ8tm+EYlcSL0LlP8qY6tpXK3JYo7C1ak6OqvcUEdzWQ57RG+FLr13fClkR2/+/qCpgdq+
1sSObPY4Ng8HEgmvkpEaEgzoabDbRQjUJqIDUXIbjYLzFSvDwUWzhBHjTeY3CV2qYzaw3Edb1TbJ
Jq6+1NnYj+kG+2Yp4UsGwE3CR7bZeS3jvZjokZe38lZx17YiRBYQtUHIW36Ra47Sr82Y8KSIRjTx
aUyOsc4W8MwuFXXPbEmdNK/azlvKtx2oYd04NHMDFvFX5iusW3USwEUVyTxpLF/41I7q+seoL3Et
5Tk2XWkpHnsmPlKp/43eSP0Oi6Fpqqyjiy0Bo+Z8FvfV+sglQZ+FU1dNkBXqMC/uXjHHKfqLyWDL
YSHIUQbK/DlHOoG0/p+FaDALM0TI0XYPaYdye2xwXij9XyW7EsWR9wwkxua4a569Na1CAkccBR4h
ly9yAwXhY2RNnJyEC2cW5b5Pix/a3Bz8MTTD454JqU6bm4wV8EZ0CdxImBpfEOqNXshinxK/Qe5l
VoKsWtX98zJ/P2WI9FqpQebm9XF/7hcL9a0Wj/1mhDuljQQJYUezrzXaaHnw4mPxswjPz+cxyQf0
6lVw61xgLUIoiSd2GyzOsNV9bssL1klTNpuWsKWCHeYlXJkheaXJ0wx5Z9/mkXXU7z/tVszB184n
zG4931SvIlH0xZYoPUDwyEZ3G3+8K6r24Uq09o4jAdXTY+GyBv1IPyDjZAwIHWpqtn8FZJ/JLlQu
8sXCo3OQmXumeBbX9td117/PqFjt/Spq+xWER7bYtM/D9bD4LJ3Y810rDYt8sZPF/1m17AH/6tkR
adSpQ4NQvyGMC11S15W6dxVQiBcU5XnOCekb902M6rv0OnljBj8/O5X9HwkNvCVZRzPVi6E5S7Da
LIlrf3tYZUvR7iwO/z/DNeuhrEEDu2PfI1PdaeRUQ9z9MJowtI8zDibfRFS5XZW1/TIKjhwxxBZY
aU59woeCIyqZQyfH+r0RuOOATRmUGhEs1sEVLGk2Aay3lkBAkY1UHpIiTLqfZwaPZp+EflucLoE7
izdPuv4c00R6bb+rJnlyuZep6vny9krIGh4fWDFST2k6B1ODxHJ5f8HTT0sqPetUBCVLfYR0NOtX
tSHbwgKIVGcaa6cUApkpNDuhxoBwL8QMIPxJRXaXt/hThZHZFCeFdYa9D8u62mGn3e6j4C+1IhFU
pJ1dquWkNFquXLNd0gMzwAIhxU7f2GDlgeLbh9EyFUZqt4sN7cyWdWvZPKYqnmN3ITxCP1g+bXdL
4cP2oYZb0HlOwJb7sUxt/GoIfe6UKMpEQEJzHSWTlkCGV1/yH0HYS1Mo55E1MyUQtRY4kSmkfIgB
yFnaNGC3Z0d/QOSlxkoAOf72PO/acjdYoua7WLD2mLu3NLE9tZnelkMILGGUmyz66z+s4kCzK6qu
qyveyWJmckddCkF4CaMDlTvd+6hGdR0p8k/OZEMUJacSdNzYrOTJbt3K0F2x5KccYmwoKukSFK0D
xBOmUkzVUoGKy+ug3AcGcimsZf+rVajY2MaedhyAmcMikG7aVacUvqrkeSE1Rm0533yb9SdcVHL2
RJlehk5Tj/lUDPUEDnmdIqb+yRN5SjEkK/zAanqEEV4EVMr+iwKS9P6FkgcDSMdr9yn6i3ZAfOre
KlYc9/tFpIrzQKsaDEOTIAsf0bGBewEPaH5YjYs4VBX1d23uRMjkzO3irU9xeasqtaAe7LPEgHAW
td2epND9Q1wWcE6QYaLiaG69HdFURhFh65oWxe7z9oDOw15eLnlDO1OAXjXkOZbaXcPls550bi3p
mKHtSmHN1FWODnTIAB56ccZmT/awUnuSAq/pgZ5GxNxUHe819+UAk+LiyU+E2/Q6Kc3OeG/bvntR
ceWo4pZICrrXk8MqTgGRsB3q3SU/DrsCpl+0taQA7C1vI71QUFFr5zlTyEJb6UaavmENa7U16CUR
VYYeEZhmP1KVXRfosade2sz8dDl+t6zPVMgGt+BtGrB2RQ/SXLzA/zxdZJ8hvmGLtjVDJUjqxMNd
I8T85grO6qby/ACSd32Lt9Wjy1cQNDZZlWF2OBAvNs3QKZH5L2wGHTfq6gSaoGevNQK3Exez3TEC
UU8w4rp5vPUs0J+qgOaswtxWJkQrjfXJQ7mJ6JG16963GV1AVplqWsVZV2vLEiLQDdHBt9dxIxgd
SKSUYWJjTgMmDO2rzfSv4M3W6+87fi+1IU8YygEhFiXKuAqSiKSMZfoxxCZKbVyRnY32XKkiIAyk
7iXyHDJkTFlx5i7D/gwDvc4+nFlQ68k/ytfaadsEP4Q3cwpWVgAxOXDtZIP2KwY7htvBoAyzsqB6
CGLh0SM5V/ATUiODgrX5Dz0Kx7Q1WwXguiiQCo/MTDrwtrpN/XOBkIBysrauIb94V5eJLYuJ/FOS
AluxRSrC3MPPSSehYX+tu0Ti331Jhe3npl70DQ/HraZTtMLannwsnwcyxrS+qWcwZVht9ZNHAdTs
/eL37zrcg+DNDy7zyDaM+lrffPEKsHAoKUXgarSdpEQ7Al7VetwWriL9vohOU5PIE5rlTOkIccVE
xC5xgTKHGlr+3wQFh0yZVdRmH68lWR/LLBaZwn4hI0lI2GLaMB3VHiHoHITLGm9BZfxmd3eqAZ4/
Pt4ZGE7yVJObZSPzBS/JAUVQbQq3tqKRlwRtqfgyte0Ll6iU6jcWTrdF5Y05vgvzid+95mpwi959
1pEsV3vHmOan7Ag0rLtcDxWsnmtsuMvgfASK//SVB7FpFfbzkccSZrAGK68KwapnRFiP0DDw4IVZ
or17Rumet4ASkff+A7UfR5T9etU2ux0PxzUMdgY28D9V9MAbOmBUWTXRWkdwA2BDNK09MHM6WU9f
6xI5cuU6ShdEPSoh03ShSZ2AC7tVZmepr5OuLsOhjnFavf2Vy88y4YqvIKgtGbeiCDnzWoKwTr/W
aBVut+vfcJHa1m2/E6npKUPo6ai5Yc5L2AJsdZjuCRbQm1jIUQuj6G9Iv6F3QzqagK/0BQWBeWzV
RX+N4u1a2gxka6BGl9rGNO8BowkPIWKfrJPwA8GYmn9Ulj6fka5m30hWxFCVGj9DsDkvPr04hFnt
cgnpRLZKdStljv5HhR1ERQBIrZN+HZU4D9KHf5ECDSHXHP6bYik8EBagPqVHdLehLfU3Rpr4Fsms
TrvNtFV2mAQvQ/oIC11R0FpOtz6eaM56BLCtAfbfYp67qxu8hb+F2Mya//tFfOKic//eCInukfjE
epShBpms0rIMMSP2w+YtNkwMCMItuCm87g9hyFMQJPGUbtfwy2CwwdobA/G/PrR/he6HujVsVsQx
I+oreXPc0qt533cMW46IFk+uk1esn+1KwaM/ghGBMMn+EtykYjSm91cHDH8MyALThTDNoyj2O9et
hpY5u+P060+vPeNMAz/9BU/yC5ZXqLSKSEt64v3I3pegZnn4yI0giZvqsHpBavKl/ymPxRnvqQfo
T+p/k8dSu9CpxknV72Gm9gyBVptPfm9TgUfhFeImqCdzW82YczDqYQQ3C70HirjEiivNIJxYc6k2
zcyTNU/xNA9XsPcsvzDaWrJotHTaX2maGohKhIy09aZy5oQir5DkOyJNnxmmzyBXvGluHY8Z91AC
LvUaKI08VbG1tp0oNW4lS+0iH5ABXDDbE/n/PXbN8Jn9HgM9rRIUN2XnyJb6m170P/NyfTjQQjIQ
2+5Jxmwcg53b+XliU4/Mkv1c2N0qtwNT506pe3HI8WQPaYS/6TkejbZdeTNJ64jfftlxyNJcUxHn
9Om+HUmg8LAC5MU85L/F35Dyol8ALTh3xMQTJt9Zzb52xSQ6oqo2/wkmAZDkiNnr/16KMG1iEnPf
mrTy/9zLvW5fCO+abXnaLpp2IZ1D7YKSxKIQla1rQelVZ/o3KFedHZxtAkWuD0/x04NeEWeVg0cW
onsmw0NMlblBXdrxZTA2/ec9WidugTq5Ez1iWkvno25l25VDC4UO1CU1pmV0vuRtdFQ/1ZskOUjI
RU+WHaYn/eDbpmIwvpK2H4t5uXm4v0nO3c0LKp1LN35Zle2mno/TEw5O6ANxJbqbHCPGi7pmm06l
nEp042k45ZQ7ILcUsIpZG/rii75sgWNBT9lEETwRx5GWNg17Jyx04kxlmN2ztCRK7mukN7cqMQDG
6HqmjJlGwvrVHT2YLj+SsfkOy1llqsti47VqrbK/Pj9SsGusonf2+wOsLUt+7tKiiQkm9VKOOi6Q
joDSdTepdcjk9CfBSiGXrp0W+3FoMXy1a3M6BdRNhP04H1YG8NZRX4fXiioO5+aElyvcLJdfp1TL
O8DWAdCeM3g6X/9BauprnSiKwtMRi+eBeGrhRe5AbCmCCQXRRjDCjyAzz3xj9OZydZYAOUXm9mXT
KAoak3HTJal7PEbiAO3UVz4p/+EDQMwW9p5QSwdTqTJPcAzmiWyXv+BZ5Ib8UupY/9xreB095DVv
IFIqSbnUNG/0HuCKzyGkkTcivC5B9aOPspiDTsz9d4f0yll8RK4RBY/ea/nlx9wz1OVT09459paZ
c4xfDEK8nEg0mtCKond5wNKSLmEeSdbJMLG5mvtdVlwE+znZEGgXuB749dhAHniV/Ksd2v1CB6Lq
PSwNl3ex0TeVnTQCUSVSAbrcI2Z2WBD0DmmymedyQX1flYZJvL/qO2fxEuFCNu/Fn1biawSYBH7C
xmCa9qPL2LcL9vbaANqcQrWordcMUTsflTj71YhMXhdipHlIFmhX5Ezo1ztBJgZBVK7toYFGRarq
T3hVdQIXx5X+kHTuopzKHFYgd94pDCpKV5Gl9BWnaKNiFM44iCKSsx+riiH2vI5RCYGO7TS8BlnT
6NhNpkEvujUQwReXCoZaQxl963CFJezlhP9WrNQpFLd7l8pIFVucAAS/NuR8wN4g7fad5ipUzVPe
1ZGLh7rdPZqtDMaGQ7Za7otyuke3dAHiITd9O+gzPEhiFtt7jb2u3yrPcuZiYF6fcVH615w9Zmi7
y4Z/B92ScNU7zdzdO6ckkBp3G9RIUjz9V0rzFHvc1JXmmAdYnaiH00mvJ3pW1wpehgnF1JSpyTpw
nKDbwLWxmWJZS4i1Ic0DL5HyDA/0/CpTPDOvclwkTXwDBxbzO4UmikUYk77vmIACTfJN7ZxXBYQr
nblvqV/0Yw1saDVPiWRLq7VOD3QtBsHVgZCEdNPIdvM6lbSBFjqK9RUU8f1wR9KAiivBJ1ftbzFq
d5RUEMfVM6YP2UujLMuO0w7GtGuDW/D3HzQfEcARoPvv3k3hlo9+lNow99Sl6z5fGjXPm556STK3
gQ/maW+jNRijSYCQulYs6+P4xE65BqcTXWe8rmZtW03aJjvCV3ZkspBMkwXO2/uIQmqcSDlL++K5
RiAuXbFRsFtFpyyRQ0mJgOaB5fQOM8ps4vyZ5lR9ZiW6bjsTX57DcbS3zQoaP4qZSF9N9iq89o9+
rOwt/ry0cug1naKXAsa9FZb1m3IPERvhVFwA6KXlSOCND/fXydSEVxbUjZaQHkAZZtwy0hEYL34V
COyGa1QLatjoLXkH3k/StTH3HLFugU77dx941A13tOtau6dBE3zWvtN+IVH3d4KxxOnfxojhH8G9
LhDe7rnQPzDDMCF3zFFb5NWPQVCWYqVBpF9IDbxkzOfyHRUOaBafqJMKDzEZNQ3NyRopK2gyImgc
WlrT05K7QPEpE9rvuhAtsW5wyjspjMeovO6dkA/vjXBpqmBApmIhyI5g42iqvtD7Gk2rEILwymkA
YdRbUW9l6Y1xKK7kKAkCJAaXhqpsBYs0zhuK1SMweWvFHtK6tTPkNVYdu7DboU/mk9eGmMy75nlp
yMCWlwI/8t+8PINaVX5W6FwjSengfWpVxbPHc/YzaQF9PGthU/6lIAVxfs7/HmDT1SRyOwMZJF1h
avz2XM/3C83kUfiB3c1jaWKk9HZtyOE98hlZ5nzXPGEkmOxYL2TgzyIlSwEbMmScjEpuA1SqoRUR
VTuKekP8jaGuwCVcyK6a1Fj+76NtKyomqU0iQ0hGA/aDD5o2usJ7LhzZd0/u5bxfAB2c81wrM6wm
ifvvICiLiuYmmyvWzWgx0Clgs0TplV5eehql7NefQq2H0uj9RXvt+/WsFPRw2XTTSw05xOKZNKeU
iqfrCewOlE9WzKJEw51kyuLxx6GljHXXpw27Fr0VA/ij9syIgC6MoBss6aPjo54LiQ4RuveLNbIj
YdkEmeDHoL/76jeviHGcAmCjNJp9ASD22Ieil6PmgLfGghduHV9cjG+Px0QVlMETuzYQnzsEsqav
LD0wnA9QPm9bn3U2AA5r5daHA/kK/ZFBJM9O/DDwIgTvmtYuTNh7jgQ7q0bBgqyXCIKwu+aym60+
IDRDcXVQl1R99ijPdeGNH4kWxsUSxxIiMqTwgiIzm4JTJG7TPc/zIVrUS84MP0M5O7k6PmFU4eYq
gddzqxhDiVsxLN98/RsqU8kqebspLOQza8Z8e0qYwHEZYRo03EoNNDIy++tpfmhgVaC2cOK9wmhg
auDu76YIFcGtgKD2/THj/te3fT8p5c9FJ1GNB+VAVaDXett+rD2IZ5ZHu7p1DNCNE/GMv8DguKQd
Xw7s826d5M40O58uNF5Hh4yxcBUBTvDaOz46O0Tqe5F7/O1PqvqexQXPsElJt1j8CMuhRZrjvDOB
K/Uv+kaA681d60IRGqQ2jiiLKAIs/bfTxD3EaOxf5Xt9LV5ckS9UbhbnZtvhmAcjdcsmXyHpS73Y
5YpaDXoziEjRZh/CfadkQ2hBnPYOKgEUWGsDG9dPN9+L/fj8b8n+7YY79K/gOIC15+SiIC2MYiQD
ybkhuMW8z3cVRJZCruYE6g2GtNRlphUY+ci/p5uD6yJwJME3qCFOzPhDzToLYtV/We/dBfu22aI5
SpT5fsVVnq3pcjLHm9q9O3yQoQaAKBcDxCbwE6+lExIKkO3DAQuD9qfY/QF3NyUqxeUNVsxHQ+nl
/sDqavXvLdCfEe83zMrdU2S3YwlswA+o8Nbu+lr20gjfsmWLHGSG8qjs3w7jNt/IE3Z7m4TTB3N2
dIrmJHa8lFK4D38M8CFXwMrimpVUD+MxF3I0EkjrTL8YM2KdbLmxqZdKQkZjHRv5G8gR8Oc2H1OL
WzrVJCvZP9X2/xEuFgBCgSqP5eq3I+aJeX6JXS2b9gDGeRjExwOTyCG7MJVP51mQ51aebgRfnLy3
dzIZdPfi4xEPi5rdO8gnMlECTX+VZNQ55TAZcrU9tAX7SZ8VBT5904r1e1CrwXq6/9NwZNs9M1cV
T97H7VwK7oedkYwF8dD6onQNPOnjb9y41wz14cB8Z5J4HEcf39zhYwrHAJaiFbOoYk3lWg7HI/vb
8AGNLgp0toTDpg2R95kVv1N4akVCn/9VHaR7EbNuTxU0MKKuzXBrFF4A93Pde2hmVvKD8wmebJG7
3Fw1h5fNiKYUyjVDEf9QPy3ldHFp4kQ2x8i7337nsPOer9ZoBx8K2xurY7j0Wklb8I+ijPEpEvby
n7WwYsm4BFhdbe+dQ+UMjllhZEIVr5uXAsSBqx0zJZv9sfqv5hCths9b48iBmP6g2N9sRwR1e4sp
W3u3LcjcvTMFAr4FdEMlbZe8Q2BAPtVTytQ4EkOwM9Q6H8SBuR9edSDq7lWnHJ4l07mdxUf33hkV
AphYCVNHPzPPseOPzkgDjkZTEim88YJwZFLx25ZooRD/OyKKSbhc6KQfTVjzwKCdPd4C+ruWlNiS
oXBzE5Gu0HshxwLoaxroRIi97rUeD4dP5JxDHOVJel8K6kaFx79xRUHb+QmMWP1zGAuiHUKcBmHR
RYM9muVavB6Js2oakyqt9g3YgkbQdKybBbVW34Y9QFqFPoTk2nB1dMMGxuPvkX7FL00B9Jtz1GIn
yqE6sQ/xuwiGibKTa8kSh7gicpvt4RpgmYycRENt59r4iiDlC1hUMZWp2zsKx5Hfb97UoLAkPi9+
ttoLP8ipuE+xdf9c/raOQtZ1Lbdv196JWwINbdPowq8n/ICHiIe59DhSual3ylO/oP+EJ/4M+aR/
BCvzmSxQnRZCuk/MzBbA4It1/b51v0q+PeoOvDTZMevh18ZI0ohR9sCEtasiwPurw57uLfmsGbWc
Pr4C9UmTy5l7xSuWwZZBPJhjuP4lnF8YWRiGvirBNWUxkVbz+RQyD14zRB0e0IvghENxvQ2+zMhc
lPuDwB0CkVqEb9x3Q/wJzZByNEaAUn9iQ1qvk8tC1okwLYg+EZjQhBRmbGgg8AiTucoTT2bPPtw8
eLVFcrdOGvLtvwYkG82kgTG3ctWZWKpx0RlNqyi6bsnzKa8RT7DG00ymcObHWASxH4kdOTKEHhNb
FshbpQp2t9ebXvg7cIPVDoxEw/njQL8UPinRrluTL9ikFd4Lqhva46xQw7wghxCDdM8OosR1b/q5
KsbZGvHx8WtK66gEu7r5ZkkOmLRk8FkzpYC8zSpR2UWCYMLRdMnAJ6sz49SQlgmI7HmPZ5pAbcj1
WI2L6VI/gilMb87W/jn+4BuW4ftViT67uB/FIkg8f8gWUqdzh3XvYJVNXVswH82rhxhMUH+c2819
VtfdqhZPr56ptienzVSU0rEFqHrYeogOcDBTaLczZZPFDXG88fRqXxpl1nTsOnhbxDCMnZ9qXSaX
sXbaMZCO3gtyA/fVBnIBdVZJZ84LtHRiFqmhPFWTku7T5JzojfoOnaP9u+H4LNzvQeFN4SKQ3BbM
v9DkDG5sNoGfz6PMXu7YLKyTP7rSTtj+21MfEbxx/8xdEp2Kn1eLhgzFOhNvfrYFVKRUt5c4sWlB
6VZ9Rowo/NkWE45SsxK7Hsd/NM1amK0Fgcwa9aXce6ei6Ei1wXJ5QLzALHV49Dqn+z/Tribo43eg
RdL3a+WJXQeAdSoHTQiekWjqJUK4Uek2425+/du7uzTagMXqP5v+av30tiNVmXO5CQe7F/AJz6tO
vfsW2OtiBYLkyRZInJbILmKKfigzaRW+qRxX+xiY+E4bhuvRZVxp7dpH2N6Q/8hmFzcHlWiNDoL4
FTld4lCOqY5PVq5xnSGnXrlJiSvIGVkymmM2yVEMi85WDIOhJuktON12CiRB3r9FdpTKmUKfDAlr
Wlm5Vbytd1uX8si0C4OBH6lQuKKtO4dtPkjruAeO5tPau6VOznI57J1h3yHt9Mx+RSPV8fPyd3IQ
iXTA6eZhqG5GYwfA/ytLT5KkU8gRbFOuLtPOedXGfhZ5UByeNrt7Y+c8ul12kVPsh+mRcmF7HaWT
k4yZ0F8aWWAVgRo/mIqs/yjRlIwNcYn4b5MPyjhD3TQttuFJYNilCd3BMYxo23DMBqvqkz+pPN2u
eFEkkHLODZEHVjKiuwOVELcp+YtYXZcuP9InmVo6pNxKlaJQfNbt9eRM0WwOnZXI+/pKDdrWCsit
CJBTnZPIcQGeWIVqBAjDphljcmoJSUbheatTlYnTW6Y7Vk4PWGzHPp5UM+QhicvcvdMnDa2T9H9G
M6RZ2C2VJYlc1YNKV5fXtWoRoHALAhTB49pIE0rRwdawp0+yoKCwxT5STYQ2fKKYkq5b8RYFeVbT
GmxwaQx9RiBhkQ/3sMVx/IBfer80j0IjTY7SdX7Rn4bvIXZbmyTx/Khs0a7h2uKTiBNVcZBufcZh
d9uct+j5+8f48DhwEVyqX17gIROgaRcbTZ/ESw9lBjJGMirYsWz2CgVSEKKTtZI+CXbRewmslgBo
Ql5/l1j4ywBVvPQltK5eowFxFIyO8456/npxOlWFBL050kqPfJ4YJB16kLFb4evz4gWHSlzGbLmQ
2vVpzPaxJv1kl9//PQBzT/2EUDgU7EmDp3g0q4C6vP96IZPKCB0Yla8jdhNfOEslJmIu/ZU2ft2t
IPdEuaB6WxtRjcYX06okzdQ5JfbD0AxfQat7RLxOcrBs246grNaAxaW3ZE4J6gNrjiIauqrP++RS
+zfKPlyi29OTNCj37fvj0fyxdXlfOOwrgI7CqcoGrfjzOZtjt9pjBnl4jMLp1xxPrIeItaWJubPp
BMDJKf0wnpCErc38qNjy176s0u6AlmejlTRBT+xHv54KEY0WenqdBeRl2RS6PLHcQbIz2jm71P7H
Xwt9VCxJIbXkdO5X1D1vLeqV+70a1x6Wjp+r6I86FpdKu/EEJmrJYR2NhExwob/oUdGfaQSxJYEo
6u3GlnjEA69+vf7a3M2lLKnSxnEDQm9l0bfTIpx+Mqtng613qggT7gPeY/MG2dX/j67I2qTmpvGb
bnuP9U+NJpoURVSV3KPN8RtW71chK2QFb5DMjItBbAEd9H29gRlH5Dn+oiB6e8PUpm5XDcUStsOU
X3hBBRcqB/o6V1t7rT3oI5fixDA+pj7KJnC4RisKfddLrsyOfQmhqqnp8JuriUjMk+SzBO3udooX
Px65ndaZ5kjIrmDhbZh/3mR96Nm1f1TSZHxJaKtok/p+rnEtnP2zI9CRFd+N4VmrmMCI4fTXcuPu
bKUItT4pF4TSZwgDjrPxCd78S8Rd9k/7y2fHsoY/7FfCUoJq/kMSj3pybLCDORy1rhcYiJQKp2LW
/6OnSbHJmmOqoJQ5LHoF36AIc1RA3+Q0ig/Kcy2nv77dvQiDvwNSXx5a+N7IXOuEb7KgJnvAAX3U
JjMxxFgagoLgNARvBVi699t03PIoXQap+STkjpP5ufCGiCrMr2CMC8BYkhWTzchi6UfQ7MTUOQoD
kcEY4ibZ50b3GGMtFq3HuWY2kQJhUaQPkCz4V99tkBe6wqdX6fST6ZQq2El5t3ka7TRS9cNdUn8L
a5b5ZPu08skjiMtkuvNjGH0WSbpvzxy/djxfiaT+cwhTeZKfYeihr2veKQwWsIYhjwxirBNegUrz
sM9d8EEnq5Jc/bUOKjIN90jvonL0/ULisxRy/trvltTDVIdaIgK9oQH/z3Q2cssOiVVqx/ByKdFc
iMF/ieMnqbpB1gyDz98mi5ZgYkzScD0Ji5x8wfaGLjqZupfn0ENfAh8m8ATii62AfLR6va/JwXBn
RZCSQF2nAS81h5nCwzmS3oRgxrWXB4R8qqHLWFzqun1+u3k5y3QiyeTO3+QSc5IcAf+sApK1sZtT
RtGE7lN7pBMLE5vcmgmIz1zlvweureW7beQNxeS6sxZBAkXAlbvuhmIy5LraK1t8FlJnQb5Qj4lU
xUOme27fibeYLpizXK8tIUUXDySVt6ZPgR3ngzWAG842DuELWcs67+JIgwMm5EGb6Acb+UW25Q0o
HnFpowXfXS5wX3jQ6VDHxc9mz9H6QyhLFfXTH4Fg0IKEefKSIgJBfHZIZHhPOjy6nKat3ontu1xK
+bMBxVRVrlO7Y+7F6w/57WWv5sUdQb0mI9BuXgjYS2AdoInTXj6ivpuMs0SzAvvotNn1bZH8Hpcd
Ik/SWUn6jurHDP1dC8Fn8UQQHogCSloMtsAXvUUcSQQQ4U0cfobX28zXJMdI06sL+lRqsf1+YPcP
Wi8HGiJuolMVxSzy0pfST84PtWULYZSI4JY1WZ35bPoi7WjcPwmBP+LNY6gd1lIyPyNn1RUJhtN1
aOsifOzGNqJwFZfQrzzbykBnHGxjf/8V1cuhPR4goYimfYNMppGVg774o6b6AXoSMi+kDA2eq2kU
kz5BlRK2lnExOHl434uqUjfrHUmgzkBMgvaHfILW1+T1VOZyXAFovr7iAtonPTgZXhHWYKI/QF4h
1TdHa8pvPG9fyPnAkmDdUjPGRpHgJ0fZriIQuN8krwpucqnOWSvgU1KDP1+iiGOjNfcbQ15XMMpJ
9x498tp3YyHQ2lZt6Emq/+2f/vbwgZBW1I8soV/C7EgmIPJmC/dOs299lb+s3GmVHsFLOJBbpzKe
sm/iaLRuMKrfDlI8IwHd7iouOcLzt4bpNavlI2WilWP7Bn1gcAlqGENzsqHlbOBeguE09KJQeZ61
+D/8+1PsSfSKmJUdYmWBBpKxqjmuVGFKj1/cssWtuTW509cEESSdkiScpeUfCcLwrKstntYvYje8
ey6NtjwV03uQ7Gv9Zg4wFBlfLTlE3HUYWI3UI1VKeNUFuGfUwYdG2YokL/piYOtbpWY4J9oCxL5k
SsTJj0eq2bd92Vfb9Sq1abXEvgDa+BuYu5S13IMHw18FhcU8s5uM0cQhEasRP0Rc9nWFfl578W5o
IPuyAwjxeJFRfBC03u61hI7Vt7OUGdX3+3xAt7YFzPKBJssIKEbye9qIoKRG4+XYndxwKA1Oirri
b2W9Ait0EVugj+ywXLBNXAx5Y1i6qE4rk+ZeeZxA2czRVv9YQyNGgVqZhdh7+d1wOwFD+iBcgmZR
6v6Oq+BgqVRtlmDzL1bfIFfsSa/eodLezFEr+uA4ARVrYTGp3yz68NoVtLptj+ip8fh8mM7KChMs
+AOgJuqAv/Yw+w8LvU67eBzDs6o63WcoeR8bJ8857X6/SEeJ4V1jndVSTqcKuWJnpqatc/1kxvWD
2ucMZFhM+ULs7PLCsK9F00M+VRPkiyED9Jj3OBp+ou3fRSU8mQ6oV7YCAinBYQ2j+5InSeDxBGgc
BlFmkQi1FjyZFhAy6I2KEkN9YpASVc9lO18YAoSARS0gpCTGzGOqVTuhj6B1CtX8/n0hLH/pRjXS
ke9TAF98V4DztltDpdP6LDkvJcPsCxXstfK1PPBSthnz4j53vkow/s1XaB0vKiz8RjyfzoFLl29T
GCBNfU23qAT+wmyOVIKXBiKTZukiaOcLUZDJkukz+P0C7rYvmLr9kuzNnZQmD49PzEnFi0GQDwCJ
wUooKj2ROEA6h12+tWjblpHb3qH/tFjEeJWWxj18aE6JldTUtKoYSrRc4E9jOi7twi+GApqY4oCm
OlQ3WV1BOXqkf3bmX6r/eVmKgRs+/dNWhVKnykcqC3Zv9I87CPAqXuj6FCrTm7V4atz0Zg+3pam/
Slhz3SN6vbc23VWS/zh0bV+xdcVci8jg5JXNt5rhS5BGdCNZSIRImPTd1IUOHG64JA3GDVl62pXQ
E6wiH0Qn/Yj3HHGEMgQTCP4CF++FvvqOt+TI5S08SfEU9b3SzAUDNzDTvXlatvsSyrPJ6qTgEIyS
EfZj3NzPqoxfHn7Tc/OSU+ztB2AwLm3n1hAzjSG+71f2qMXW3qSlT61qLjd5mdw01dMB7AWjNQVY
gJVJh1yX/3h1AFOOuuHEeMwjVQy5Y0WDswxQsrG3iI41z3PxEc+Ow58RiuKtx15W7viZWsedMkEU
JZ58NKVyUHZhiHjoeF2Yd/qGdp8JHg4I9zJDBKJBuHHrSjJYtv4viyr9r4MJfnxl2REh9+6M3Jt5
QGcdL34403C8Z024fZyYnLzMgjVITxzwSADDHxCKGKXetY8rHzSXhZ425OyQkTEwYOBkW/qwamPm
sCDvHSBHnXbbG/SWE68oGgVNxTIkoDeabrW7VAl8s7JoiNJLNxpbVEfEYGHqsPKF01ib8N0tEcEx
fT7O10JhWIwNJuWldZxrcsUP386wO8ofMafJupwICwiA6xEfH/BTBFQflum5Mbfc+/cAvT5VEIlH
y7NrYd9tpwwZmtN53IBnLaltIKQ2E7ocGnWw0Zdr4FijRUv2heevXcL6Trt4IdRANZrCjL2aTQv/
Py+zF2ueefb1HxDRg100b7N85M+pl2DNavM6Scl449cwJW40P+7dyNeBBEWoBhQcX8cvW/XOE0Rj
8aMXgrYsIV2fJ2gkVKuN3P4T1MwyRr5Mdpe3yAVidpRylzLP+YTpNs6x9nwXVNj01/ZfT8+RgQoC
NAGMCcquCyN3D6G8S4lndI+90TBSjBbVxFDcIH6Rs5q26WqXAGAxY3N9pfcOHDBjFj2DZ3ICMNbB
CoUkqfyzR/C5cpAop+3ytfKonRmlZIsJDakGn3VBjJ7AmZRjEmBbeQ3JVWuRwpIf+ftquIC6tkRY
K7bRo5jIvFP2aefHTe8bQeb9EYhbMlLrW5YEkeFz2iEhDXJSvBxL2XF0HC9qu9jXVQ0RDXzgKcn2
n3PFGZtJXNvEPVMYgXQVYGwsfIdF9reiwj2eFSV22kFVFzq1nMFCQ/ohm+uSFPEeldO4V+/HWB66
kldQ1tHhuQT0ZmQhBd29VsRcJSCZgOD2txL6GHfHfdhFkdg9SvqcUJmBZp7FAIABCfBWHqIRE+fF
R9fyETOmPmbY5uj9i1cgsuDuPy1L5nXPb+JNtPWczE/aHni2ABx3Tes1+0woWOf1CRoBj6dcjvV+
P+0TGb7jUgY2ndXaGuGyVpYWxjNiIzf/5YxROwRSACV4IKRZ/PVaIr2tLFxuGArL+iMchbgW2UxS
vQXDLNzzpInIF4ukZYonN3a+aHkGpsQ1XHLGMRMyrNQd/44a52tPHW2ZWg2dhYwFRUOvm98bPB6m
+qW4X+WaGyjP8wnJtn+6jpOyYzW/lADcwFO2LH22FQaXg0q7hJnZLMMLTbPlMG2B0lR8Eh79BunT
elegSSPZhO4IwRH7xaylztHxoL6bz3h111FsOCTLxHm6T7Tx2V4G8fVPqrBeC/5+r2bYZ4loADT7
BDGF/ypb84oVTiFPqpcTftQWJuxy3F0szlJ4wYjXSA/dC1KVk7RJA2WeNxaFeGHzjVjhpAMrsy1f
1P3v54w3bYi96U8y3gd3+I+HVz4P9Nl0MeeYOAN/fEPOl76B6Zks7D8qk2vcwsnrTKssl3BIpuZT
3FCX3OXh1c6+ELGPJViM1wKJpFht9EIWC0SZlcxj5CsBZbJnV7weY5ufVyP6dmbupSo8H1BcaopT
+Iz8aN6HZ1ng4MCez5qCKLmFxoWwz435DyHFHWV9cx/B5LGJJM/ZNoAMEE9VTj3Qi7l0k0IIpFBu
Xpc4xpUwehwBlmPeyRZVtIWA4k6wQXkb6Ixqt0Qzhd+ksUOjeaW4Z5Z1ELiMoDJ/N4yOJ2NkpE8c
8dD/n38Epnxte+jBEA6zetcroVjOGGEiW2iqJaE7tnym8irC5GY3oVRhKW527A+0yI10XcvBdtWo
buRHwZlkRVMFVc63vW6JXF/kdO3kGIwC2XbQodDj7avHxZfwtTK3jx/6DnKrXul1hpqlp9u5BMVB
rUz5weTI8qwqq5CgRDTprUbVoYHpqQg29aikSLlqC16WFaACuhVvVHEdnw00hM6IYvKepukNm885
1l7febKWBiKGvk/MRknkRDe2v1D/yLSsRx40gwkC42V4oYUz1pi6qGiGlSbiBk2OaTVwuy9rGLmV
m4FtR8pANFirHhsm61tpVurQg8vsZVXkmL8I1rKSTlx8rpWN6/Sbg0DMssWzg8CHa86tlTMGLG1f
EhQt5TJ0qnCkKfD8ZcFBnJzxFT9Kak9TxsWgtmibIEtBgCDgYvdQB+DBqeGT/H/ECIpg0/jbxmph
tLflSxg4cM7RedmCqhZp8LEE2tIcuJYnyHBaG827wDRx9AQ1w44Xk3sVtHYxynpXpN+DMGFyMfnx
gXNf0cNV7+92vCy1QYBuME84qbrOCAl5is7q2w3OWnFjSF4qrEoQlnKF+sYfZjf5WgEs/AcWcVB5
hECeLx0XUiQQc8ifIrcjdsXXpF7JrXpxC90gtmzMCfRSuYcekaiESUI0GDdDQnZrxo+X/4Zt/4Vi
TXq/m1zpSOK9ufWJgdn9pB64TwTRQQ5NPhe3/L+cwY7yTzEt+tCoHNv2ZCWhgb2arjBHh/LnIGE6
Xb0i7XqAuJe791kZ8QZaFwv3BXRPR+7euf9zcIoYDSaCTLRMbx6jq/7YaRpzaSgzzsN/TPFklRNc
e+MBfpCS8tq+qujCkpve4HkvbTqbpJkzgSBYCgg8f4jXI2NA5PO/D0OSyH4AX7kfVnf9gvZ0e8jC
iGBSMtTJnMN1bmYpcZC5yT5CNiSfUbInG7q/qJf7hXA78IHCx8q5z1zLlGMgY60IL7eKCiOKXyPQ
eroSgkZZvfcowN+2j/J/EcWorpzWiCg9B27qQqyacA+KCpQwl/M5B6lpR9oZFWm5zoxsdyAUbehn
ZrT3MfRPanKZBaSTPVB/wkQAD0Q9Q6vNnKzq2mXWTBP9127ddClnIZbtM9aoAO3gXbIco0IvqgfG
6Us2BEkepi2S0d2NfwsBh5k8dMhvDI9drBfMeY0z679SoEo2OH1tW8yr/gYi52P/6Zj1zkrNIefg
T/v1D6GRENl8HHBoaZ8sgIn71LOu7/t0Lbw14GF6Zc7AmBszXliVarCBOqFDaUPXSYI1B1arQaOh
t/NFwSejEiM95HmDtlJ2czcCJW1D0okivGlNIG47eCNPlGzw969SnQ6fJ70rnzedFOY4aV7VYMTh
bwYLv4TtbMmSVzxUq4/rcYt87QwByvCHiUQ9rLLbhcgXyISvVrMeLV8MDD6v5vAY7JKjXlPBi4m3
Xa15Qe69wN5HnywyzN4hTXOCt7+9Mqn1/eGkQ5QcNn4PSXpl9QeXGrp2NKzf0KDBOA2K6FVPrp9z
ajChjN8nrprYt3zdO4dmlG/DKYiF+cU8g440h8SIvO4+49/SdL3JUJ8193UFwVbzBZDUl6nvSkEo
9HjQgTX9ZJOr1L1CDdlBwS7AksSLETPD/1RM3m8DZq5LWsgf21Gbyj9d3/iTNIhMHtPnfYNp24TN
G5P1lOGOPm6RtfoVgaqj8LYoV9yicHK2BPybcpkYza0zNmbW1VESK9irPqZ++QHTMl9iZYcaEZp9
SFIxbpIPE/LN2UgrO9d3/acQPYfCwPOoIMTNxY8SS8IMSuJ6K6mc3k1zm0joOBTo7gQHuXJ7s0e0
mx/GYZlDkKPWhgQimh5JDYDdkHvAZuhYghkNb7S12LNC4PMSLsqBYRzboSlvRNuUvmjk2DNYVl6L
RHHAlYdYNlxXpS6Tvz5A/IsN+NYIJ/j18cRImnQc/Ej0R/exT5pR1iIdjKlDRg4XjXJQ7l56AuzF
4UZ2oZRvraRX6HAQF/Nf3JWKze2vzqBiMglfGvEz01C2WcGcQGpFogpKrQi7TqWUHmUoJr1mIbo8
+eoumIzVWMV1HHm2xccBuGp6bBK2yW78LaNT2iwtvS5BomZhWt7pZm2G+4bFWwBaSy9QNVBgFRSe
f3nfFkMFt5gkvTb771rn5blIKTtNE03m3cRwmY2/xyOki7JpjN9il8ZeOoQDECZDYYrLxNmiSTVX
RfV63FyEM1EEKibAHs/Hpo7DsGhpxo7goEkQ/3ZkqYlQrtVh2e0BxJCF0Saf9YM5sxjTXnHnlbtg
hHVGjgj0TOPoqffspf+czOFaB/A7tvoBVUylrS23lx1Pozu5H1Yozf6Q3wcTRShae0it+NJuAQ23
eiCXxe3C8zIhdfZ8pwrCzaHMsx1p1VurffSc/fmFLCwM/qlV5w6BsEebOZK1zgPNfWgSZ62fOh4x
rxxPsAanZkl5+LHkljxGu0trwZfkUZjQsI1s22/qoX6P8cwhtmdpz0/F/kUORYiGr1iutXY6Ib3p
Sr90bDLOeR0DyOsTn2P4R5oOBpaqSgfj+gDmrtRiyu2A0ZjzW4lls5z9f6v/N6E6j977ItwKvl9O
7vR3B4GsWWdZJ7qXDn0l+j3mEEbvZkYDwO3rOsJ3XBaGF2SVAQ+3CdzmxAkm5hVBCcUQe+1M2bH3
mzVyO5wXs769/wO76o+FYF/Gz1R5EBWUHAZo1DkF4yjPdGCqu00qW/Dojg/oh640Dq30ziBCS9wQ
TubnrrmWqrpTGATsJIi7Y8CmGdLpZtOdNpnax7RDqbz9xWI+AgKASzSjVmN40IiM7e4FC2AKRW8L
747e9lBYPQKEJf4vfGA+qoyYDkCdmvpqynu/JG/FRs5HZoOxa0agfZl3m0ynt+uUPbT8udv0CIns
zfKYsVmW9bxMSgqHUSp5rqvnn2xE4o/CxzaV8pbs6TmVGuGa5K7nfYhUX/zrhAhad3bA+VS6W9lP
bldcihxA0e4b8JZulUtBvck4fXXh2oK9ink/Z2Ctfc7pmBjU/WzGlgn+pAMs6IR18JIAGZAaakM5
0OO6izKV+clqn/+wDEMwl3oxj+hBkb0sWL4puEu6Tgyx0jv+fo+gu2XoclNghu38UDgCci6PgDYT
Q6NjGA+ACLJRyRhKGwJtM3+8P9BucYdc1RGiNGXkv3HLgF1TZCSypmIbYxRGmvzguEANjad1o1ML
JNkuuNaScHTzT4Gy5OIUkxQjX2TmE7s33nhEzrc8lj+uW/M+7vejJNXmpyx4mu37gENv4M4N2X3y
6P6ejDHifjPGTLH8kWfAo9kWM5ey9VGtSVw/ZNnZMY+oeqmrotCO5Wj4pH9XS+3eDIQuAtBmgF58
wqv0CzBo2LjcdY5Z5Dpnjv4vjJlGsUfnn4vl+JsVFIB7FUqtJR/9mCSdefFX8v+TTlifYoiniTKY
zZ6HuC+ZWLu/ktKpwznWmOUs3N67CCiunQ+sNUFbczkmVnGKSkPICrAJTkbRfQVteZKIwTnqWAxj
0oZROzGYHCfb2+zCate7+GrHZUAV8DzBfAhiNWvIqYRzbx+yw0Nmllb8C7xbgHUV//V4ECHR+iQ/
+bZglZzLon3pcggt7k8hU1BSDhYKGhhDVZqpYojd7BlNWQESbuUHAOzpqPlUaVrIZVS3u9uuKAzQ
vOAgssM244fKyrWfOCac77jyQDrBN9o6VDr/n2xsYczpDU+9ub+agztO6Vdlpx0UpdxdEapzHq9Z
wZHiqGGQl2Opi+KT6IK9Vr3YyvlAwa8qv9WXFHIr5XR0D53iUqAoT49ubLdcojO5w+O24Teew4Bf
rIKxneG1wjo7rBd75aQf9ldhrbmD6J/lL0wajzWKvzlkK3lUSJPf89v9Xhb73wRc/TEDLfxko9CH
N7m/n91pTvFH37GR9y45pjbreA401VUeCeb5oyZuSC+6jMctcGo4QSk9h3S9mShv/mqGiW1aIVZp
KOmFpC/tjHDykNvzhy5RYx7ZC0N43v+TRf2ByupAtXA/oO3bnesGK7w2v9nJ2ijDO/XqZB+y6LI5
SrT9FyfOEnSMcQEr3TDRiCdrxhLdtaNXGKUIcelSwB3snYL0Oj/DNwVCS6jNFBIUliveBAJI3gYT
OznNN8nvmrBrCLzwPuuFoRtVuouIoylCzO0LERpFxd4U8gxeigb++LCyo+1AYQs/O/sk0wAWN5ZH
Qyjfk1+mbfcsUKu0a60CGiiRvm/B6P/kW+k/53nvktVnUREcspxjAOZ5dPk1qMVq3eAs6KDvuf7z
kaI0c9OFBKdQY3CLAcoyRx/v+aWlxCzLvgMZamnVEJApwnVDKa2gGU9gM7gzaHLhDd6oyj2VmkVX
uHpegM1rjYEa7OlyZdC02yigmGF4KNoXbw/BvuxztVQ/mtzQGubf5cfvSKqroMBW4OJATNzhLf2g
tcyCCvJnw5XF3BvgfOro+DZphWW8K0jesFHbHokDqjacNC0/PK6ToADX75Cf6P3i8T4AmIHaNB4g
w3g3xfWoTd7VDWx8JdI/zH/Q3gHXqxNa/akFHw1D2W6cVOA3B0bi9tKR5zNF3AM6VFijRxhx7Kkt
pRSl2dyWrqSQziZXcrn/As8mUPgfBSDnOHqpX7oZwTsRztNVVW5NxHtu5yRxJCyGgE17gq2mJvaJ
atViORpOefUbalvt2Y/rIWnZ70PWJDnlNjuFVoxsD5Z9+XKKqE+rW6t8BDFR7VMSgHVekEAsqI/v
zIOjAlMvdGN6Sf8wUd5+5zio2zoc9sKvXjbnzXyoZUpW/JGxrmNVx/6pL9hWyeY9ZSza6vjymz4M
sOig2lpVlieQaqxpODNSOZ4sdaacgyI+we1cQDI7DirHsOjkO8T7Qnb/OgbxVx4jwTL7bOqa0t2E
z7xEUcnwu+6AvuC0p7SOf9Wqn0GyU+NwyYM9togfgdHULiSMa0i9XYpOWLi5qvnZgzvBs+nUctkn
3irXdWZD31cRZdWncb71gnOAqFIlHEIEXTB4OgmDSDXgWeBF3HC7Zl8hqTcdVVlgA8rfGryc1aWU
EefK0wfUctq2m2DvZc/RwhOT9cEVb/RqbxqKK+PWy4jdFpOO1+ZwVa/mCkTc/XGX0/R8WrZ7O0FK
XrIyW7U7QcNRiXu/JSLHHfRN0yNyvLV1fEauG65TY4KSIIwklmiRvI6EgNrBWi2he+9OMybqkKkQ
qHjZ923dsyiCV3DuIpgnCvfRPbvEKEvggkB6zQrrA3hpWsVvvAfZj84biW3kq9AuzuX6iCcex6OL
ujLLM+BQiTODd4Jcl2FhhUN9VBJtFlYmm+X08tnegoHaKsglyajH6akUWtOi5Z3jW4Ve465htzUE
5MAB1Khi9y75zkWOVgROKchyf3JpDlHDseQBF4rBDShWn4vquspvldXKmC9/0YgMM4/qyft065Ib
FL8n/04EIZR+03W/Au2gVpGcLmD3u0/MgjL3V3b/aTEOtbBAkLwvZL+v+w3xUT5JgUfi0ubi+8yq
BJ93wFLaXq9f6haYauv1Ju791dWXFpcl1gWhqL/aSktsEBkD58RoES3T5EjutzqkzJ9pm23+fpME
M32Ye/lW1iADnmpvcp26HVz0rPgz4Ds8V2e3Ws4O4tinhLxBc6IzfGuqcSVLz3aOGR3GW6sFHf/F
KqcEAOLsVtyENO5nuvYHsErLJsw+9bS538wmczfLtRzQIArHqZUXqhOs+eSrbZNubxR4h1MxR/TS
VKR6bJ5U0+dGMyhL362Yematnsr04p/n2evVwzT37SY6zB/QIKRBE85xcmGZX/dq9y7fqUwcIe7x
JZlY59JUJ3YPjnpTa4jyD+jyuVQcx4ZisFh7iX9/QDLm+c6n3aIEgr/K6WNVH1uJ+WlWP9MOgUtJ
oT4Gn3eb10H3qx1iS0tiHsvxtERp5l6PLCva8jn9VNSsBlwUwm6LOqi98DNAQWZR174VnG0GUESw
J9Y1U4DbCDtCcY+w5c6A+DORlB48DHUMYoF+XLzmNcJfrRcYn5lzor6yxpIlwpYT4NMSTooDBfxC
dSad8nAEQ2/53LCsY1vX3hmCAFkIf0rjjOlZ4eKvs7tjJ1RF96VqXeT2LKcSdVElabneGHfsLFet
kJcj5Hec7HLugCPgXYyLDJ+j4347cfLhajUmUEbOULR0Touu+6WUNuhDfWy1o0rmNnO9JeovHjFS
lNVyeDLXHsrZceJOIBGAoP8dso1bwX8bx8OC5Doxl14BcJ8fqsULuzSqF9Ie6LTCHzzV1qKMa0bC
PEfl45rfDCLlGr4h4BNjsdZXyZrHWqgCWojnXrnn/6Va9qFOicS5NAJ+mxDuwjLzEzfXVdwJ3c6N
hDDt19GMCNanmabj3yEzDv6TQCzWL8FS3QPWYmgEfIfw7fwlBeLHI1/U+Y5lP7FB4VwJB64Qf3WJ
35fGbNtk6u1k6rowGTYi6RMtK0a+eLM1TbbUQJzY28LrS+GJ50TH2IK+DfFyf4kqmAkr5wjqr+NO
7Y5Tv/tCCFqtjE4HX4XXb9G1yK+SEDLx0sgYTvCKr8atvDEly5XpnSs/RYH5F7tkZQ5giTIysIcx
EA46uTe7rXErDEPk/s2aIhBE0ZV8Uw8Kf0320iASxbh65Rjws8fyAcsfWlVfIja1hOjYXA7wUvk5
3LhUN+aHcRhfuFauXm2RkLosUckS6pUuCyBh0aAWicM3MmJYQlMXazwrJNiHy77kNROmtjoZxs40
B5WpnT1GxYlwf1vXDrNBfJMiBoY0lyiAPfrtjzRdEiK2Veu6yv7kxqwEq7KEUtZey5+flu18Y0HL
hnkZ10bXMaikei3CXDAMcoRHn2hOvl4Afz7GBTHrP09I++wpu1H0kR0lsa+li8lkvw5ckkNn8EDc
YnZGDk366NEgf1ktP8cu7C0+40IwUnQKxzT9xYGkok8IdrIDMawutvxU5ywZA+bRtL2tIYn86htq
GCwFN92fr9bxlcpNrJv6pYaLyIxnzF1/cpzqOm3/5/mG6qpPuEdwM1f4xKu5A5pRCGTAOSJtV5xV
IcNjFJwtm6muuHql7CxA90oJ1qhp4laJiI4rs+KbN+FroEgzUZKdkqtbJgrkwzOk9N8LAfCncqu1
Dd47g7JC692h2ug0QrkCEzcEU+tbvqXfRcEFbsfE7/Zp0lWfAqt56sWaow6XqFtjhTXv39bzLb1Y
++v/YTlcJEjHXy1rM+isycZBTFa7sgokfH7eJxDzWvth4JhjGHGkZ9uR6l/pso5VQSnVdy/4x8AU
5lmzpLRBXA7X5KWue8OV974pBr+FuZkUySieNHzMmBf65FL3Vd0MR8imJkClEmu5U+bHQqnjV8x4
kFja/S95bBfbkmM87YIqABk7SnrxKNoNAl5AjhOjTTtIZmm/TG30MNGH6FLsZhEwrLAOWV1FOsS3
huLVbMYzsVgUAC5aOyXuzfO4i5KgIqm4GB4g8To+XxhkVjr1drsasN2/xgNsVwG5aA8ZmgBuRsSe
zZtAUKZ17iksBOFQu0VQ+MN4vf9Lw9Y5C9kk3mD7RogvShWXhcahG1mEHgbtWQpdwfek9IjkQKew
XXaheCmEtQ+N2NH9jHr/qTqvm+jS90AN3C82JGH3m70NJyHL1W0DhnRYySvtnyIwI2qZ8/uAHUkH
Z7eDkiYbmuQb7R5wX29rI/YX4igsROVfqtV1YEKZtsDAbCvffH+bdwFMpcaggjERmsXm6iYXq75t
3jl15Km/IGl65PFDwHYAEjYdI4V/FPb3oMGFX9H6fOOLY5AhVGHLOj5tCLVa6BlbxRn4Y9N/v//l
MUwWaCI6sXxpACDtYkQiy/QatuugKoSH2r4zdmN1T0YFK/3WYzXszxJX8l00LazsHgdv3AUFqiqR
J5pULb5itC2dLMYCIQ3uM9vW6xhMZnH/QalPlQ8Ko+0+XIJVlM8MnwytNDLcTTZ8Ki3rmG7L+KDF
Qm3h73p/pOziq88uF4AUlseICl/t1Dj5GQzs8C6eZddjEvPZV7T6FUEJp+Is4pDd3aEBkQIN1R35
55JqPdihTvGa0Kx8sMTjNpuH8QftHChSHJ3nHs4YIJGzIDsHErUXt2BsQJlmWq94yRvUSSA74xsy
90sOmZuMObJ8cm0QJHlOxFdj5xfYkrf1ejVtofwRj1a9KFNzAchT7hdhyJwEX2JHKGKv+dQqzfB5
hfSzQSti5orX7sxNGd36QrweqPvdw7vZxotsLmuB6nR0VX1AOiOqnGrSaLdfjY6UG9/UA+KF/RAi
fMO6tbmUWFKCnr+0TWfjmE+8xXDu9Lmwg4ZB2mjS07ASVqjJDO0my5XNKdfKhmitF7J1lqnqashC
4ZY+nu55I5HOsUOroA+bIc6c46ApTjMkAlDbqhp/evZQTf1LQMso3d/bNY0eit9GKHEjr343Tap7
Om3hPcByu3lV+Pf1/MtLhs8wvXjZP/0vSaNYL4mstHILq7aPfhKsTvFH+GXCR7rF4mTVt+3VBVMW
Tg36a5M3OGmT7ZABKeCIpTt9gj0mwiLEQ5qBPaxELW94Pc+pMl0EQH7FG+R7FNgRspX4s+TLSJSm
MvJiYcmgrCWTGmerQNYSBA/WrQC/R0w0jAFXwmeIVpm2SsJp+7+/gbI7e5p5mXhMVy9ZK0/clWa4
YPMHzMmz+0IurrwKPhI4aCYYB2h09DGTFNQe1EvZMbxsPy4odGh6hLwgsQ5aqwmC8Vt0lAibPV1u
HEy/a5Y9MsrgqJ8KiNADmeDFIUDE1xM7hlNNYsr1vmbucgOutE7AIW11yaqof6j7lgDLSoIVRKR8
YEoQ/pwadlY39YpZA+lz4gmC+7HyAkM+adrWnqO3BwJggtBPqwZOrf77P5yfoiMhqctaj9mmJZmZ
k2l5kCgvVtEYUGZYfch/jCc3wN/SvXXZ6XtyqYoRC9+BYBkpON1KueKdRYubPlnfVg0IunsS0j0h
aUgleYtfuoFAD3JsHKi7v7wxPbIPs3mi1PC6z2XVttA0TVvesXQzttnhDMFkG32Xj3TbRy8VWnra
+rFNHNXb8uOHjZp7p7Y+Ne18zGD980ZK8ETQMDXCiepiLTNZCvtH+hyi9XC3UjGqE9SvEvrt/trU
uZHlN13vwyP4OORXAXCU4VPjmYgAukuZGVyse1CTclmp2gr4Cx5dHzHbU5MWG5Sx1lZeB5NL9ldf
GTtXpuY4EFeIwNtN868ZYFipnhh60yBkugWbLoap4B9JiZk1AX5EdD6372H9jGZeJ09nam9xyE8n
bwNkXcxExpXB0ZF4/K0gPNygLvZ24XivayjJYrdTGZySgN3MPfQodlVJuVTxXiSXj+eBeHe24PLU
DT6aJSCybstZFjC5mYWQghZszkcTZ/jyaM9/Mlmc/YIm2H3Dyx/ne3irr4xpHImYErkkd/o6aH1p
MZHnqqKPyo3ROBIxLK3jKhGnHEBkm6xIG5oJz2FnyGJnOtoL0WqulWQ3kjFUIPSbByYnsOCl0IHB
ej34jOCiED+jw/pAdQcMuwsyIFY4aP+Ma6dgxHO+1J7zUGs15qlnmRtKW1IRng4KFPqdee0lfmRb
9E0Qr9gUu9gmc9dIRRfGZBsqWXjYh5b16JFhrYPx8K72GvxJzMicjoyBAdQ+jI0Z0EeF0QYNeRfQ
SzbPiTB/y8d/O1DR57yGuJ98JDz07yqilGLjHmvNOD2weLBjORytz6x1qUqsCGhirR9zdFCNdgZN
MuJJZe61g2z6mWmjMWmxg4HcuPe56meQMWvd+bcezMHwzMfsQz8wIHbcpFscvaztQZLs6iFPZyQw
jvEDvHWvRDitowkKINw/6ZmkRG4MA8sPjdxReGVK4QkilI4sIiFs9bGK7bkNn9jHZJXmBjlvJwQq
Bse5YCGYGqe3gz4HfaOHUXxfh0JsmMtwF7uh86UQt6TT8ow6mM5QR5SfyJkMaoyZSbWtnxH6JQHt
T2YI+D8k+ySaGUBVzzkTrw1zQhez1MK7MRs9TDWf3P489PFbjPvjvxf6E/Kgy5bCLbytE2kkn2Eu
ZniK0FlLOtEVBzIG22o4dBgnHdN8fTRLcw4LB8sH+NSkdfghBYjdcu4ESTZ4Xnu7GOsSKNp93G8n
+g2XwTmQTdOet+XIqDpnQTAi9DCKVAWqjI2Xcu7iHu4KLd8WzUmtFRZwTj79lhX42PnH3p6IXnai
wxijOzb2T4LMuk+mszBXymkIPjmfUTLeZPojkhZUbnrMLKzlCfvJFNpcZSzfHlg+HN/L0yV4x3zX
/d+uJwpzKu/RJOSRNsJeiiCtswZO+wdwAfU6fnl+g30G2EUf4swdS4yNquau++KLi2I68U+LIVrx
ROIKkgjNR1ifqpfsMspYIJEjqrYDaaR1c6zJc7pf3JkK8SNt7235P5vVMxSlwyQf83+3/aq8lkSd
WBgu6cPZznN00glfu83JbSzOXvMwG7WBBatLco5ZzkqL0gqK/I16ie8nhPLDrXMweHIJ3iGXtMp+
1rKKZtAZZzJ8UgNue5sNiD6YI/XgD/RBiQopLzGSEJX6YkUC/9784zbbxVDSH39/Cglb6q7TbmaT
xgjtqclMLV194Vj5RgeixYNVUhfSqhRW3ED32rBcLyoSD5DlT5ytbBGpkQpFN3I4v8PTwm9sqCR8
jn0Fa0oAMkcTOxU8aCSfgrdnbPGHd5BnpOgGj8iqEZ4uXuWnt4eZwRjgJiH5J9hNiW8/nh5pJN4b
PQ11CeZDxuw+thWL/p9FcHrA6XPV+tp+WLCSDR/zx5i0dSvQoniBFMhSnl4syslLAEeaaMeIi5Zm
W1M+3/oFfQwyPOgRuRKmEfYgfUvYw69jA0RQgv6WoAp7jQCnzuGlXHZ5JzKtiWBHcRJq1I5ONl30
lm6p840C6FXe+al83kIyfRmO2lNhhQOxH1u5jtB0tPmzeq/ij1PcBhpWnE8b2c4U4mio/dzYeiIe
t3hDVWvU37nzJmIHNRpv4crk4KszOzBvBW63dSMJBWVirzlA0e2VBayOSxh/0lkCJqY5xDXOdOyH
yDMkPf5FCH4UEcvlPfXHCX8VT0yBLtElm14QKFV729A/vXLQvaYUQwyUwUJ9y+VtrLNCneqeKbsc
nYFLh1jmGaxpD+tsMQ+22LCJmCbCuW5+5U7f1EuSBuXQ6LAdeKl116puVtxi0pbCrv+Mb3GlZYv+
z4qLiu2irFQSOU/s2G+0M7K9Ppz/GqOMOKNMBYnk794YZL16ECyc0pkXK7HkBDg7e3ra3rBIVRV8
+9aooVzcpRMH5E8m0QDTp2xQIDa0G945/cCi+/BE+6K1liBYmu3SJ6hx+AJ/wK5u1ItZATC3tvut
JeOL6XMKzihjj3TtimqHVGtS8MgPPeuLlXtoswH9ROTpVGvSTghYL12wlHB38JeL5pMoy04poHJW
5nGgXAPuGDF3hP/XX09gNJO6lo7t4P/JWMk/94cv6Jg5o9+zvfpPFsN+LDLkoA/oWGsgbQb9N8wy
On0fZvN1qZzRFVxMm9UzFRIyIaKoE3UqF+VtFTt8CTBjuz5UgTdivdbOUIZXang+Gv/NSPNwZK9N
ejFCJcV8wr6MHpazut20xdkXrFPdWdeK0rcPSRqvhDtO/zocKBlu9pqOeFFWobuLHfwq/1sQKk9a
x2kIGjdDFosSjdzPcf6J3SXYBBTb1J4vSzrOrptb0QRc4U5JT6JrxWP3qBpDRnZu9myvJ2RKEy5W
1eet0Ws1GdZBCOoQpREV+ND3OkBv5UuiTxKjoKBP6fhJ5kVG3/0aCYf8IpBlD37IIN8W9pNyCtEs
zFqjRw+Gb7+99ujh4jAeIoQlDLv5LIf4j7z2obgHJ9Ztqa6QzHOT8cMX+RFvfnjI27hBK6Wf/8Jx
MTOsYmU3Z+tzg/XVMwpmPSAZAtO0eOj3mKudPhUQX6oT4qeQ/ew+K176CNWCcXP60yC9RwuakU7K
MgupdS5uuO872yzF9YxKYJg2Rcg0DOhfZRWYLLpWaDLvIQfJ1ZAM3l4UQXB10Pc/qfHWGJ6vQ7kR
E2zVKpesGJWoG8FnCLQFTumTybTfYj14mbinUisCsrOFSWegJ9A2eUG6DyMYtLoAyVraqlfxBVXS
vfoQ3K/YgwFzChcaEzhvcKOPQq0jIExBtFIec2jEVyGt8J3b9dAVJ7jyxGmjYWNL9l4lNcuGPpQS
umqoIwSM/gMld/yKeGsF+C6JQxypWzJjwq/jo0dfRvxEVwVrbWfn1zrnAtPPlJVeIx/g9/OryLJZ
zin1Qf+yFkmm3cMOVfZSqqa262QedYJN3wFlIJ8836uDszpMkHRpUqxQ333vSYRytYjVK/HzJqH+
QxmkiuNePKPAqNHCk3sIHBgEcNAyZVuN0R11JvwhYOFY3jn24fx5ADbQ/u3QV9gySxV4/H1nRZKj
hdW1fB6Dt+6kIXAeYvhQZFyytMpIt1kycXn3Tbs0I9jMAb77Bi5Y1V6kuF3yevWdwGLPwiYgh/xF
AJiFxGnpH0E3cpUri34ZJkMBkb61Q+K+9YznOeJY316MWYXa2mQghUGwmMXzqIIqZrDlqZxsEkuN
moSkPbUMeHqlFPBI4/ehNpFRp3hKNF16FGuUuB8++k+Q0f6eBzcZgw1DiJ0DykWk76CE6lkqoRsZ
CX80tJfTQfEd2e1k0p9fYHxOOYcqUrgyhyTMp3IzIEFjV9N9TdVAiaAV27aQ4eE4sGpaOc968ZIe
8El3GuWRUvHobxxSp4LkNYl+jzwei2juGUUZ1b7sHuHLhZFXloj/a96pVPQpAJfnxU6rEkydMzMA
FJapG99UzxjQEP+9QIuXbbpqn80fU8nh5hr4n4Al2hxViBo6jOc1bMJvQrChf7eFMLIMWpwJ3e7+
S9WpAZyvhXMCgLL37Kbnf4fDG2pxySximAisAka7ENPJo6P5Ff7Rr9UZjHUCp8UgmsJbWD1W/7PT
9b96aO6TD8QFAoFmiIUasuKLWcJAl1mrX4dVEZM7Vwad/qLqJ95KImktUPG/co5h5rZsMaBOEFzo
Ge5lsN/4slZFoVeNvO8HQv/5Lsr7aVZHkA51pm2r6Saq2ButrIxyuopayqedXR7OFx/BWych+L8m
0p2CsX5wLfzQIuqC1EbHU5Arbk7+VytKUdujKIQlqncVC3iZDBiOkFOEpoO5FscSsn67+A3xwSG8
XJBaNJAHul51oQs8fehPK70agvD8tPLYjK6KMDJ8zHdDiY46tAbikxtAVWtfBWEjRkqHszH9PvFU
Wv7/1vG9GOgDKBGBT8p6of6hGjdPmYSW47b7eHjwynN7jHnJXKQlAolCK7Gtriwyno3mpWdjQqyw
QzXlmYtMqKXflsFXrF4EP3IuX48ONXwdvd03qLP9imk+o3f2YGtt3wkTzOAK1Rj+GNlsqyNmKYuY
AyL5CF3ZYuy8NXlpdbGKWJk+llJfwq2MpviVEbCuE0ZarY5sCXTvFVm9taeAnIzlHWBCdBDuzNG/
8dfEhhf/1lTSAnzi2A+51P9gYauOjZPdIWYmZ3EGvcrIsWLkUyZj5CTpu+vnPacZZyas1XOZNzaQ
ycG/OUsn9hyYiMeu6C1mhpsBCPMftwWjHhSZGCQ8C6Y+PgeWKspLCCuXoAQprxmGeZLK/B9BcMVE
TjMOX+9Lu9AdVZOroHes1DIAXXJvVprJJIQdIFTgTxgLg4oC9A1LTiJxrdxkKH9XUhELhQVaUHMb
qhtHSFwegYDefQ1Kf+czSY1Bwf2t4LzwDp8PswwzNgpLXFdg4OQ07JxNSXtf/2l1bugsJPrcpz5v
FAWg3wBnvvdxSI9EbD1RiU7ViM4EfqljbtwaJOoixXEeHJgQ43w2MUQbv/Wa1+aRZ1lcdMCcUDXG
kamzWxYebw6Rj2tx/S7ph7NgZFL0Xh+iRscMvhvSAOzMsBlsTMigl1BfX4QH6vvqaa8h9AOat6hm
XMNSZMNVPGy6FPES5O1X8UThvsc8QFwbf7mlP+FjdMo9Bc2M1C8YKvD7Cs/au1M/p4+61N/SPTe3
1VK7y+Fl+GPWxF3LC+ulQd60lkEJ4V+qhdk+Iwh8VJ3rLKgqy51NFPOuO5/wqywBmnJHumFK1bua
3XQgUW6PeiAHHcp/PHidQuNwN0RP8Lyi86pYOpc4v/AsvqsYf26cP5MQwut0WgVBU5RN8vOa76/l
2EyjdSQdYWtBtr4uOVFpjdtGIiE/jwxOdsL4hBX0erWg65HnNLwPsAuTZfbb933rXEiHK1lBtzI9
zkzHlhaKUOu64iq8o992+4h5Iwica7tA2uch7mnphC8+HGhtNBiwfaPQuzUZh0oqD/dI/D17LJeP
ilTlPZfZgEiWpfsew/ybdpLqVRa3RFZ4w1zGl8HE7LGy10QUM8N2rWCQ4dM7mxm/axUGO0p7znGD
Msm1bQD2MJlTrks4tmu8ScH4Wbr23KbMs46hJXtEdG2/YOn86tuMftl0BwD9W2JFQcoquZDYYLGT
6vAp5HBPpYMNB7+wgP2saiQnmWjl51n1Oq60DLWsipY9Hfjw/A2upge+rDaOQtk9SMuF95mXGmW6
A2I1WMPhx4M1RdMnOuL0HtnGaRD7I6zSmhkT5olbOKwSyoqjtKXG1wwJyTcgSEo4Idg8ZacRtWjs
1zYU2WgTNUaviR1AHq4Ch9bJ9hAAw79/X7GH/ukoIe4oYFJNwfm5uNS6DgKJsC2gK3pqjIkTYTcr
lhfnM7+TBJKFCZuwp2Xi56T6bydBAEKcmLIN2Ed/dPhJbSXnEEKn1ppdhid8hU7HBUPiXB1VTVXT
PIV6b/iOIura5K8+yMvVultw8Gb8EY7K4bnjmwrh6+wQH4dqWv1WLUcuV1put668LSJMKBDBeY+Y
Hl+bvHjow1EyzikfrvhpAXJh53BJUoh7Meiup7Ib/4wbOymjSnSxZBr3FQTIkvzVHLnEhuVTR2jG
bT8EKO/sSnrM6EiWCMDrGiC277Aw0N/49IhuuEJOe3n7cq77IM0uBr3L57T2WJO2IngNiz0hF1kb
+KGKvmU4U3tl9GQ4Mn+Y/pco5aktqr7y0zp8ug5MGlUlg/PhROyytdIUCVT/z3GEtIy/uPTXijnd
OtimbBWJztJ5ustvBPTxotGb2+xUn7rH2YQAfdovmos3Z0SswW70BvwCMHI8fZWhVt/TV64nHPVn
zka9T/t2rcPPM0v+wH4igDcxHYOyMPS3mBD9SRV8ZVPuGG747NcV49SfSrZ+2sCmOpB459elZF5P
aqCGWkOcjtBaOFRTW7l3c16zlXPy/5z/o1JTl/D2KjEBsQv4Rk1uO65obxMXEkoKjp4t/8pjGqfE
d00NVZkijRwUV16VMwaRARTiKygTBArotBPNlWVQYkWd+ybsKaj4sy/56xOHjkgyJIZAHUjzydNh
1GhpA7NSy0PdxSdUDgedNWhyHb6R9G2Dw6cGvu+owmjxxTuImHlOmhwbvWjo7VfsXFCsEcd7TAX7
fNqUr5fz5kvqliEpQ496hHefj16vDXF/XABLqlIKABBivWHzyRy9/vNyq660/RK+YBcR+6UrDM29
CK+UzVXJf3KyTa54dDO0+hIlV4WVmHnzJaaphFKQX4WqOIFzKbdPHRXNv77c90Y5mcPXbXAE1jhW
tC6HqFCpwuQKV3K58/sq4wC52RdwCApTWCH3WIud5bpYwAHH/LfFjOiG41PxX5nRz+Z0p0UaETxC
VPkt02SbyjtVE4MD8J9MJIUEkBrCSLNX1rhse3qzmWw6YXsKe4bqT+A9Q1esL3q+c+ETIpEezWup
E+NOxOHp+pJK5X21fVkUGQeDuu18QgWmf1n+KBtSnjn+1ev4m+Zh5se8oyxDLbvS5Ap4TpMh0MW9
7glJTUE3uerBYPSmO7Ukn8x/MAQZgRTlRLrRZiYoz+tABVdUSP8Np3RnYFSS/PTDzPGaJMTvnNaL
dkk7qc43c1xAznVXGlzK/xOHVz/JPfUHqkILbUQIatYEVoY113lFj0wevH4GAO/TrdjmG1KKtVHg
d1izYZw3B/UK5CwAVWQt8QAV2JesikDvxR/KgBbXZ3IaEnSOsihkRI4AVLFgLbpb5p/iOtCAT/l+
qyu4s2sJxf1NYnNasDvqNw83tsj2aqj2jNfdWwvClEALTpo+L3IovV4HJQTZGltOWhYf+ovnOZL7
pkYJd0y9d0WozaNMeRfwVZ1D9RrqJhdSUZonEIp8yBvaiz6auytPSCcdm8dbaVJyIlRrfRW8dM7E
rHweyp4sP1ft/heYhUh3+6jHljlwQKnNdOHT0VY8bNv+uhSnZ+gXxDy0SA63cs9ZyswgYZ6MHOGd
BXYKQE/SSuKEIW11aAR207joO/G6sw7fZmG7NuhcmPnH2UjgF5A0JoXQKj/95W2wxrWuWb4Or9m2
ashFt8UWngK95bXUbkr0uUatMSdLK/OP++sPB1WcQZnHzFJaCL2FmJBHY0tZfpzBZ37+3PjJGG0q
KgFMl3RQVOO8wpL3a/qxo/vKw/JFIKY9N7knHlIIqqh8QLHEfiNSfoKwkZB+ueveQO0jaICAxkT+
KfOyI26h3rYGnErrzPpKl1fIGjNutRASvhD5S7gQsynGACoutceLhPdjeaGA/zsBf6VI9pZY7g/W
uk+iKT3ZHyEcOt0GMSJvMBI55FqcUNIOc4vtDn4X40Ou8+YcANOd8vVF8fQ9un3RrAMyq5NjBeGQ
93KnSu82JqMhts3Wy/Drd8mWCTC9kU83rZyOjZX2v4srpogyd0tr+/AA1bGzrVe9OP9dmcHKXZMz
7eCu4jp10o4FfG6rBk7M8zYymQYF1vFUifKoaxnXhERE/xUM5NOJzPVMK5TTOcSO07sbxH6Y+MuU
dnNYC26E4ooY/LlD3O7Qvla9xK8BxQ1mPDzPLJjbBmaNQok2q4bHmNJFBT/zD1zCWTHh62pvQEZ0
figMAOaci2oYrusWj4XWpFLOBczjvbcywqyBVJETz3cjBK6UKc2N34+LfWzJU4jtHFya0kSBHJxx
i1lA6ZFVLMW8ZuW7ndA+RdiEgik5GIN8Cvr9rZaoajrtpzN/I0WNqyuUBxK/neHNm82O+Ee4hiqr
0eQIn2etOJ/H6tSKpl04aAFAxhKhEKeF+1H76ejNyPXrtMANeKdRPyEhIXeXg1DR6K+zYJSy6htf
Yw9cGKR7EJJgEXtBvKu8YlwpctEiO5YLxIBRHgd3DMjYgSuFonqH1cFs4yspC4AOOnik06/aHEqT
1PlzFGvURiJx2YM7TA/7eHX/L40RiXMvjMIcV41PuMkjhqkmyQ6StiNTSvxtFPhpp8D4an8lRgut
SDg5groR+ANKXBFK5G7Kc3Ljb+srNWv14mmaNAppTGTGy1a1r3gIwSwCv1dcDEBJ0n6kArlqeipC
dLV3NY20WyRvQ4ZcPkYpflICdnQ0bpEiCrC3NhwEBkRmxPkWEA4G6xTUas3bNjpvnlj8O36Z3UiX
vv3007jEB0+J+tCtNPaLHbWIunz7FrP5VmVm36yKQVnrpWkBRJK2ztKBaXKDguyj3wS/vVrzNq1/
v0fu/Ms32+LbHp17/TmkV50N9OQ1/FAsEtvdPH/vAq06g0oHYjl81ICgZdiiHhI5nwtPT5UUoA0P
NdfMwI60C4/977/4AD1FQbIoM8sfmRIEoC7VM3f2b8xUkQ8FPiyiUEGfmP2OZkF4wdXTXgMGvwht
Cr9zjviq4qrqxpZQmwkyiv+fpwsLrkcmBSJVaAWzrNmLhFUEn90FwNbTefU6fY0wK7kLEvlA/QH5
CQOrG6GYMmPLOtt+v/IgNk53+jBApzo6HVNoI6UEXa5oZgXGJOW/34K+vtR1t3eR4PNUd99woU54
qk34scBqPrCaACB7I34H3sVa2OQndT47eFiUiaUiDIQEiDgf1/5K3uyS6Q6GR3WtnFF/8OsyCROr
q5fCEzDvJFbAfDOCF4xm4z4etv8F7X2U1I+vjk0kFscVuv5VLR19VtDz6kr/ciITW6HcnlRMbf7P
4US1XvRd3rKndUJg02agVz+TF5GUvpvgo+4h2WUxngpdZSz6aaAUdv+nTCueQuS/5o4vrQjQoqaZ
ID9V5ccrNRZxAbX2QUxbL/08lwpFRr+a69w0wjNdHcEjY9sOsy6y3MQ8tH2M5GCTPRrRV/M+v2LK
1Hn3LeNBhJV8I373Hm06BIMAvdXef49jbkxn4Ofs0R86G1UmRbxLu+A2I+V2hOaI1PqXDlB0r1WZ
+oi8Sp7sXNZWMw13RHXsWxteWA2bOrYhbjub9hDLaI4DRKsrdwaUJKHCEXSKFI7Nor1DsxpuBRy1
RUpODhL8zlpMGqjpzrCNZOUU+Y0ST3nNlPsCosuqP9nmyyD9wdlVFI5nGSwTdBTCCWosfxZhn1vd
ytIMKbPq+7BOcayNMo2In10oIoFO9T2TpCLgiXmFlYoo23z4NiNGrmcetFVwRqiqcdWuP7/GTIQY
CqjFT7l6hm0Yd5+xjblrzuAChHTc1Gjvmk7DouRO4l9eY0FQnMBvyc0Cz6M5ETPRI9vDAylA5WCX
n8Q/1rZ7rmJBMNT/ZP5hIEdhFwoc9KZDu9Ojq2EWMXTp5FUQ6wESzU4oPWwWw1uU//gkY2VN7EYH
baOtv7634J/82HBGnXvS5Qlyk3aj4d8uW4aoesy9XuDacFJUoiedgSzkS8/BKXPpDe1sMapxVHDX
anQ8mV5+IlihesWT2ewCSK5r+VvYYHuOWJYYHeyQbWHoOZAuhnABOFFsnh4VdZU9jVe7SHtFBN6x
QO706euhmoQ4hJk9SZ8n8rB2yNLZFSd0JIuFzO94IrTSI+kzd3Y6EqQhEM3Mu/QiuWuZRLtZI3oE
zEA0SLRDdNhp6j2sdQcj0qvTJMJAVdMLdUxtxgZZV6K/OiTgFHZa49fGjJPbjADWKuZv1na6Ztd2
2JudS6iO5cUkRtzXeNuUsw4A6oo1xTGH7DHcx+qRRXTsESGYilNNacNlGpgDgYl++cN/JN5GqwOG
0lNlXttVIpqPEvHTC8EWO/eZXSRbvkfj84XGBxElbZxmUqHx7zQ2iBkqNYSDfvz+1JizQi2YBahf
wF1CAu4JRjWLFL9Eyu2KLxoNwUhqqy02jiT/FvJombRjiJLKUB/rKKTVo/17We72PK0FqJnBUQEe
m93JcvESzoGEW/BTHnnTcbvTZcLVtUVp/GExaJapzTEw+7Sn9ohjvha+MJZz8C3hupD3nhBRP/IB
gCAQaAMJTqz+mtCCvpenJSRMBaOe3WCcxmaSGrO/3R5ffFOCRK34zNp6ft+rlb1FTnrvzO4WiIfe
Mjq1WvkXYO092YwYyFqFT5TYdSQUMTCJg0CLxbchJaqQgqdkDeJttUFpiJb0r01AglueqFi5cVvz
2DFKt+jupJrHyHiA+aGIr3vHmyujcUerVkedOvNl9tGyh+BPWoNz9zyeniSxmtqLISbE+v2mJrgr
OSyJyHGEN7zW4+pPAnNQhA+dAa5XcX3e5SNUgiAmfvJt13PcAATtTBGFHAIyoDIo/Myx4P+Qh7Ym
Xgb7xMjc2NmGsPhf9R97Ym7IpBDtvYjhFpcJnx/5e95BNgTanxAigfjQHRcM5Fxg6rdv24s+p2CB
8rpPzo3bm/NQG61r1RMzqqpRKp9f5S5I5Uhq2T96qriY0WuslWugIj1bLy8hwp91Vjd0UIevhEyP
dRzTR7FJHCKd+E3FdgACSVDtJ7TpYbnY6XJrjP3oKCuoi97rqmGpTLhFE+bFd9M0DDvIWBabsSdH
/TVjilXbXwxwIXpI3s/6kunGs2WpNmZ3mTdkUCuZ8wVs4lPwnOBVUv5o/AwV5+oi0fWvoJbiyNDw
W07jHcESojRniLJbe60voUpz37iRIDzNH5rI25ndy24if5W0v1eIbV5WBDnbCE46gFqVxqx/D2Fc
hPpFi75D+HJgsb0p6r3p+F5q7vsYFRaql3Twjc0BO5SdSg/eUN6JoX5EDyBDvecLgSCD84xfREbd
V4Zi82pD8YQYFZrzzMVPB3WKSVGxjCsRP0u1Livvlfy93Vj8hJuTtqw0CqmoKbFoYg4DusBDJl3K
IQnZWW/qI2CcGFXKDrGwZ6Jnx+x4nKRVRdLZ1z3//B2RDCEbxQ5q3eKIC4dH0shKykbA+c4Vem3W
9ap6CHJJ3Td/YlparZbRXWtHvZ3G1VPIuLcbaf4cExYeSnPWCOxJfIuGYvvupKUy1KPliFDMGirx
lS1WqZ88VuzE4lCqL1Hs5n7nl+flDLuF/zORHHFCMTwJE3uXLICVGd6p+jxseKXyws6nCLyOoup/
CrJzkGPkMUZkte/F88bHsm1nTBTvgqv6PXH37GucXXTZFvv3nnc2zZc1eGK6WWehwPFCtE1zqzlx
PnIXF5v4/ThbVr6bN+nFcS+9PMRiXSVJHhbj8TFfS6qW/DFVsqAKOt792OtBEK1Q9K18dlIEGvpW
Mv6Uys6tTX8rbjvRFrrTflccIcAWD64ui995Ah6mUPc8h4thzqO0IB1NN71bXq6uU5uJ7zg17hgI
4ZDjIOO/i/vlHazuYQbyk326pSitTaEjItA/GoarIFYXYGMdx2jK7p5PEmKvHKfNHwTY+CGFa52X
iJaSN0/lvo0hp3rYHm5l61fPeUBzzpqkXKPawiOcKIycx1p0EhWqwXtpbH++2GgkOI2NyOiQ9ybZ
GbjPku1W3J48kzJSegf5fKbMwwLRn9g1fnFGKmlq82HZldRSR5VIU/Zlvo8nybVHHa0skSqlwF9I
ASYCqqJz9Zf2IpuC17T+deqhG9pY0rSu4WFO2II/mXODE7jwPBt9+sy6J7pXPgIVGcigWJ8DQ8MA
ldphVALdJyuaZdZu5YTCksT1a6HjBmc0IgCG2DtsWriYAmJqWql3U9fpxiJzKF4RBaoeyMlnENSH
QomKPpwoEREFdJ/ej2FpYi+RpKFLJku/paieD7wTHGO7YiCEeJ3pSu0AY41wDro64ayVXX2qQ7z0
sxC6NAVN861QlSdDwWitTFEg9qfVvAaJw7RIbpektYFNvyjL/LusahEwwCTKDRIQjI+jhQhJLzGE
pTh15BbDcYYh/BEJlpXjkl7NtAS17xZq/Rss2hj+MvC6HYpiZcX7sfXE/C2+Xf1w47ULuavafS+r
7ZJMX7+AseC9WQwBXt37VeUqW07Jk2qvKbsP+I8Zeph+gnEHsONut1Xac89LSAhF0Tlzyn99sNPs
Ilu+PyURVK7JbxEuJh+JEyVg/Y4cFtdoyin2lrTl5EfIS3M0kYDMDuGgijnufJ6PEc2VvzDsKpeM
lOWIdwRhPyW8w5LmZhpQIZHE3d5YJ5aTdlNck4RL6T4kbzHwzfv7JgWcvRXbqN+y04P3/wLwCCc8
Oh2XTZ6imDruVPHs+k/uwhpdyIS4NIK67WuI/p7dv/1riWM+NHZdpU3o5D8BMzTePC/1bOdElxnZ
zU/PQiv4yamZc/Y0qCBpvKDGS9VfeB1Up3yZc0PicxJPj+W+H69TqbMjrV4gfBkL9K3W0l15CJnR
3NPR59VkpjRYwz+PlAdcdcooD/Xm+MHSaeIaGVdwLQooLsXcWKD3928IezmygHdmFR4rMN0Al9vZ
Q0hdnNed2/tjhC89ZQXs0LJXtnGLdzbmjG0FLAHvEgQ/pzBs/XMiZL4mNGxJ3lDErawT2Vj7TLDm
0zIDKtAPdPF0BRN64r0vrwh3nqNCA6HrsAI3stfOa9S0FxUwAWT8rBCR0J4E3jSnKKdRJP3q0pu6
1AoyLhKByWo/X+TnDZX9SReWj8OJihwymF0QgObbeiPOdeF8qc0kqNK355tsRwLP3fTj7xZCSqmx
eY4Ip1XFYPY4+ctoiwgZ63ZE267GVTZwxg8Q6Z8/MbXuYh4R2cxEM2IX7WV20fwluOVy2Uyv6lCq
+w6ngaGKmIB/cHfcU/atLDy/OS282TpU5eha8aNyuh+YT9Frpj/AV2hkSfmaYrnwsTZ/4cPLuyn7
xrQqSPqCmzl6SwxHu2egCj2xjqz5uWW0F5lsxRdT1e3lcVQ6wCXbNDVTgILzYdrpYNNtT95RKV9N
KB7A9HoSxx2+yjSpHTTpRviHCsBoCrCAoxX5OLHHLUwxmbi0+o+UagIccFF3TzzgYR2lJp0elpLY
TLb85JyFeeNxb4tqll6OxY7f6WQcO87XYBYqVBlu144L9Y9C37/eaRDZvjqSXUTU80gS6MtqHqpw
AKSHvE2EGvPF1N2igsF49/tbftU9Xi01NkuFgH0C0nD6+MOoS57GCY1VI5BS9XDymGAlNW/XvRQi
YjsJY/oyuaHC+JpPpr8L4URQCbQp9b7cUdSBTUmtFubD+bOXSgWfZUUvRVwOn+eQijfbMHs76P+1
0Q3pmGbJB9FO+DbFgxDQBgab/zdh/NSA9vTVJfRsg0PUboknbwbGImrvCHQAKMR+EK3yi62HYkvZ
19rImzdxE3UgAPbGU00Es4F7vvr6tz2b7I28ueRXiQp7ZKOM4+on+T5EKiutJ4pNwuLArI4N2heb
zMmZFTheQZvWPv0GLGKwiHCGTwI8iNh7PEE7INNe/2brX777o3E5SClL2X1bXEfr4cfhBrdtWqlI
vQ20w4clU7evT/y9LhItDLQN9E3DMHupeEx6slPCbK4CpX/IJdiX8fmGbkNH4E4om46qDhQsTY37
nlWsIw5YM3IkzauWnjewL3Sh9cIdUXfGS4wIU2HbZG7QNtkw3KhihX3uX8TLgofGrNZVLY/6FAmf
RXn1V4zBM6mAShplQFAbdvlSkwkDo2/W++iWOGAuZq0YefCKhmjXhTNLmuFMAeEbqZrK+J5ZM+n0
uOxW4wYX7pPBQJ+cQCYqCxF5OIvAFSFxGZnghOcjzf3rQW8Nv+67VM4MwEYog0X8wzqwRDNo7tjD
oYoDhS/ehxT4B+w6lkDv7HUxvVAE2PblDFFacgNUzllj1HSj0Im1LRr6z00/yFzM49byAnzTiErU
w75pHCCBbb17ZsXLbBz9WQd3yCqZlWBtezWUc+qMCFQUDZPlXDGMT1iiVUBbnBaY35UiOYy9uYr2
clvH47dfEUYv0KnebUaXPGO2JZ7s2ytIrGfx9fnbImzjNT+PFRpG+bCSgJF5NnECbQLWMI2YJMPa
df6kW2OMU+mMlk43JnxuecMZhJ2q/X/QXPvqkZswj5Na26cX14c3aaZ177dHz9QnMGHXVx4waI5I
1Hyq+mK+xU8HQbWyBep9uDodeO0swv0lh6WsR4SMseRRN2NOulWAxVaP8Mv2tBkDB8JQ6V9EGZbh
dLL30icUbwGQ3Epc9s39h2L5DtAEqorZVC/8/ALQPeQ2FDOMBYcyvTI4c2sNwyfF9k5FYoHrR/3S
KrLfvbZsjCGK/BHNC/rA59Xnn3Odv1DHEK2am6jlYpbzgiyi6VORGhjllR/B6wCw20vCS+oI4MGx
F/6mvFVc22AMF/nxdf01jtN0NwYP8yFElseOCaABEsm0TF8S1h+YITQVAQsBcUBQ9fJfmbTY5L9T
lpL2eroyH9UCnbCrQMZEjNReE4xUB18FFfjNMPglv2nKzm+aPiiSQ0bnqcpCVU2kL2BWz/lB9ShM
+lI+uQdYa/izgVF1DRwS90A7DsDiGQoez//cQ8IFpf7rh6O5fX3Kv5zhyXOQxUfe5kqOIWN/6XEP
XM478/UTvwki5zA7FP3f9nKJncfvMad/4+X4in9Iq31A+9Kh1bl4AlaIxs5x1nAe9GfChwQG/o1T
Rvl0jI+Knpy/awbNfILocjGzcsq4KwDdAhXiu22hcOUzRSob9yQTk/od9YLPAXsj6n+G4P7PI63h
h0yhtXcOgys6Vikim5cls9kKwAMQOr1BFfleXf76XteKMf1tkzNiUFS27w9ladjC6py0HRB/wLs7
wSb/UarV20W4cmNGHU1y0pxZWMaNFDT+SPpx2h/5ftNwoIhs8n9ge/9hWS4wItjurinyPeJ4zc9K
RTMG2GKIqNrld9h6pSu4k0t+JOkWuWsvOMA74a9FYUxaMISpZ4DRwChn5VLKzqiTuMKTDArrzj6Q
WBOhXyEXi5y7hahmK+5DcOxbA8btODIe55Bek88ubI2s04NFcPPhRhMZB8J+DFo9xnebQM7Wk4Ce
09pUqZ1/mJbcWDfDACl8NNYenug+7pSOd0Z4TFgab12Qg11hZOQQ/TbPVRzK7ZKlZRmOwyBqrJcS
TX29UZ4+ah8NWhx+/WDs2w9Wk92jcCO+CgId0Uu06V8pqqzHZevKvOBo9zsLL+zS6rFU0EUOYac8
2Qsi6KO9ibJVvHjp0bRg+decZA8eXbHUXO+4DlcAtu8rS0CKKi7IM+PTKgE6jN11CFjEc8fBMmgB
J3JhgtMYKhOaV6qoWVW4WogcNIZ+qjWcSfO5hJuaX2nSLebFQc3aIkmCDzFeg+V89ZxEl1Bjy8T7
2hML7l197azM85ZlJ4qILDPVUa17cKgSmUOQaaoAEu29vJwexSheIKM8VmDE5ByzldBoEY2xtto4
tYQOtIRUyEDHP54gJkz1WHbwA2l1yqEZ0Hc1vr5hMC9YJxBg+q1eHNJ45Vepl1UbBrWMRnFvEwQs
Eq5v65W1UKfkcjpS5b2Gp14qyK3BvbPHjGuexo+UfkM6ABpotQsYOipixzVt9X168MbY1+VHHAJO
diYQCNQTRgS/gYCEUxzkJ1/jGlzZC9xJwXR/yY66rbHbkGRMi4frrBzfgAnYl2bvc2FltkfOICmO
YHQO9RQHA9vuD6Q0MGsL7f64OHk7DBJw7+BtzHIWMg+WvR59JTTO0myXVHVXI8efCtSUArXHYmX2
43ruy9bOkUcqprj+D/w9yPJi+4xIG2CuCoz1FaByOy2KAZAODPvZR7D+QRIZV9K5IbDFK0hQM7Uv
85NfFh/ZZzvqG+p/GHgo8Ajibm4MyUkZSoSUJeIAtlcXlxMk7bUkcVqcz8qNw/8bj6W5krXSEb+q
kO3zzEFROQ9vujWcK1i21fUIJAVUa4nKVQWx/XwyrPfxwumTDWlnWAHbmZl7Qq0dXv5FHh5toKR5
DoDWHrHaRpx/2BcyhcTLDI8l5H0HrHJeXpfCzozlgSrw88WYHJjPxP8WYjxVruBMM0FmVMVwEEix
lWJeRJl4L1zIRY+oLEefqtrRrySD5tC0IDkUhfDSF+TfcqRIDWqJ9N3/g9G8HjJ02xb+OWB770gO
eCVCP2rC3MTgQjaesOA1xZj1QdYiR9ZD0dLejSf8zsqh9nJN67xI5CwDpXoPZ3Vcng1FKgEAbQpb
y1qXG9etDSwaOT9iC7OQ4dxzWbVa52JUoShqEj4xB92d8zGpYX1UdU5p6bQ9aTQDn/UFd+m4pGw5
oGkSobwVmAvxb5TTk3/4M/Z8LEoakQdSvVdPCDwN35I/CJXBBR2wTcvitN6EmjSrq7k8sUdtwbzd
UJ0udXwRvPEZWu8wcW7zro2lVqH7q3Fxe/xGffErbyilxQQyVRx/XLIPsGV6hS+2ZzqZyfwQa6lN
nqlSJ1uW/PUojI9w37k5a4FUNypRbXpnVM61OjTLkh0PkOA2Sb7+bmKVjNE9gkxTGcwYjlU0WMno
sk70A6/GA5twU5AzZvZgmte5SRPpmRL22E9OOgjPGNRVJDEetCeKx7ntt+0wMA/nko6kuG49UG3C
MAYUodkMXYRIsm1PIiFJZPJxEOdd5D8emE14W2My9Fx5TNKKGnEzWO1pjiLSD7stqlKxiZkIG0ug
U8rFZgslQaEH+8IqnbY/V8Lbo36SlRbHP0hCEM61R5TbEzu8k/+h8exehwf6GlWh76hdib5KbOE0
XXC/AItYI8QMU3K28etSHEjbJ6amI+oIdlUva0eZ7BuCSQ4LLGbRjKOe/TUybJkqn3ZcWhGA6nUF
910A/3j5KWnV2vjE9dFkEYL6zcwBoq6vCuYwDSX1QDDun9yOPTUtvkULaCpa5SeY0UAkTmrgyrjd
3iJbVJbWeAWuEPUXQlrvLEDTL61+o23pc9D7qOg4sJ6FVpVDv6mIWaEcPI78ji+9QmAsmhOHZahW
2jFGL0SrQUnSHnw6Vd1L+taY4vEkIXLUfxhXRTtIvpiEKcNMroz4q/4hQbOqVbwmijPaULQgfFAU
R0sbFE182Abx4ljEJ2oWL14e5xCUbN+CyviPySrGouU+/lk/NS3rruhMHdmPc9lHjfgpIxT061dq
5pNcyc1TcEn+/npt4abSoTlN+tA7j4FjOte7qQJpO+VbEIHb5qbn97whKHvrTi7U1EAMVosJTlon
IUWSuK7lvG4XQbHg/LnMcHEJjNHzrBPlnIdGPxVNgt64jYsYOvan+VXphqKopBOQxqWZ7rqa1bCw
itJ5L83NcDOHEw5SxY+Z7wmhmqL+1lIX1tDVmTcnBrEZXbzLPU5dAUN+aHfOvLy/Fh8jsDxacrau
IIFLkvgW9i5Te4P1riiP9TSA1JU69S+SmUyrWojzd4C1s7t85Lm+N0ALv9jZmn+x8YZtR2MlsDCW
tUKtW+ADQC9XCMYALrTSc9P9pz5XY1XxgZPGKNvP7iUMQdCb9zalHV6GYqlc9MdiJDDI7VdOO2xa
Se0798+04Sd4BOWlgbO4cepnTcB0rT7kjjx2oJulYVV9/D/E5oHfFd7ru/a3UCHN7lEi3wASH8Z/
EIqym1qCvGq9AVs1338Sk+iThS06uU19qpLRtImbRdzXWhJGrQsbfK8vf9OB1Kgw6XwOGQMvnN5c
/8hKqDXJtKDOUjl0/s5TO28zY10N4kFVH+bcnURdYdV+WCeQUdWH6j1FzKxoJmSJAfcXHS2dNf9v
edKxzctv8GIIUu17RjYA/u1ox49pe73gM4qFjpdyCf4RB6kehPrKZcPTJMVOIhQDbRYFbRiRH4zQ
r8lDwpukdxnHtsaa6fSuvXUxewX3unR+ygyzr4x6pRamtEl0zQ1ifypotGUKJ0nh/vI1FUMa567X
lZoOLNmR8gYvlge7GwxhNPrILGQfJAJc2yBtbJNs3euePvhDWR+VJsgC33vTfXnYC77dvsDgrPKG
JW05rOQBIgf1Tevr2WvENlWECv2Kn3METSj2wUKkducmvPcWyK/gPoX+OF2wwdU9otqE8lY8ut3d
1rDyx7EnP9dRNpK6eTuGe49WPm8ZnLujQ38lchChk7hZM7BGHGweZsm2vNZKVTthM8M3N7pvbwWN
C7ZWeUeVpc3cXQxif9cf8kIuXYlcTvlj53ZBqSjKRdgYkJUhmhIggXt2NiYnUKBk2qF1dGmEdgfp
byEwDH3Awm2Yos46iAejyxgRhVDWWGkLNTvphR+TbVx9k8Jm9JC8fULqQSW/KHA5efPBzCdm9+e6
5RB8GTrSLXE5u0oq6DElFufYcQ5UR90qJ+69Z5ioan0pfzgDqUcyspkjX21kNcSbjk2mXQI1YtHJ
rJqv2piqBlW0rm/Rafy0GGJjyAs2UM82Hth26e+cMRK1z4DMDaucBKErhQVUbKCIDtOtCQJUPETf
pwkwrmHH3DmqHpg2bG2UqgGdFwCyOu3L//E5ZTad0yEFxNfvaFx5fMs9FQN8IxDjGYmop11/mk+X
fzCNIwfzf73uF1j6hFRbQx9ObOQq1H9gEZsN7jlvUGYR8GmYetRivthMUapj+MtV576oHxd+Iuy/
brrzO9Ckx9YhJCDt8E4JdR+NGktFecb1e38u9R6UEFW3nhG2NOr6xcrInqYzxyVCpBfjWL41L8b1
pQF7yAOvLM2Z2bYGD4zG0MXhKecrBbA77L32NI2yD+NAqKmQ0JGNry+XYXHv6fk34mCWs5e6jCTO
W6W8fwnSbpk1YGCUj2OYDjP2Wujcx7MX0EGuBoByQDHw/M/6VIXik2cpqdzyasGrZfaQ1rwG4nA0
NmoC28FSQ9nNWAEDT1hlHcHKfCf1J76N6dAg8aUTw4TagrEW81Eed3hsp7LGn+Z3MWDDkfpoLDDF
PLQV2NNOS5XzvWSJUhHmUm0sBuRoKJJR6Svf+kSuIebSNbe3jSy84ktXhO2JSJXvRaFeay++4ljR
LMeJGt6MkK4C8xGQZZ1NJhoH28pPOs8ydMwCf1QofDhiMcShTcxgYocie++7eEV9Y89/rb4wjjiM
zbuJDcsQQPcdAePGIe9breGgs6QrV1F+5KwbfNnlOOfGnIJRV+v/Pqr/xmGJi8xnIYQyaWj+Tz0y
zd+9GOLvNZZUDysL+0cWU3CkFlc/suloH54OCXZDjiJnHd4+pzXf9vrOMJk06212Ievc6ConRFOR
ZYo9M9HEh6KIATnn/ab3UXh5xL1I7YcqtxDZ/mpMIOVout0/8oQSYGKl4EssbQgvx/ibGHbeqmP1
2uIHIbQQgWFbQ8wXRqocqQtxIAcbTSr6aLKt3nQ/YFwR/dGXmKbqPwEZHzLJ+7VCCFWhVUymJV85
KssnPLX8xy5M/bRBCAjk7LPFJcgvKF24o5b0L84Htkv0JfeGjJCf3coTatTwBt7aS9Itmjln9PPv
uHpyq9peeq1C8qoMJu6h8wmtqVq23L5KCbpr/D/4bgiJ27XyB5PwVW3YDIKZ6RAu3yjpnjdUpYun
xTO/OU3kr+ctzo1n1G0ObcEY42he1730VYF+AfsuCo9AVyLg6MY927CFbQbu7956BG7/e8ct05Wj
W29Sp+9xo9lSisKSBEeX2LHcYanLrF57frfNW1GKmLkXDtG58kOYQdM/9RS6M3yIsqceREZKTQ/Q
LRib5tHQsaBs0XWFBx1GH4qu6ARa89NsAW6Td0rhh9h/gTG2FmVu86y6EB4++Pq+OSmgsgBHsYeg
U078U9MuSLfRlsPhsFrmk8TsmRy+DA5zU9NVefEVYZOQGVuBIGMeh1PXRi3v6dY1KN7BnTNybn/y
IS2+EMhY+aZw+tXY+25R5H8+ZMMdTnaxGbYxaNWOzdEmdyromo/zKXKuIKXvG/hXM0vFQG2ZbVih
L+d5EYVYwUcSb+dL+Ai/KKrmNR9+nsSftZP2lRU+9LTtWKd4mi45+2IIsi3HpwDPH2/MoTiv5on1
wFaxRmOw9Gfyplzq/FvknfYHq0gOkUzn5KQbQX88v7orXddGDV8bj5XsmVLMrBr//MnpzjTy4K4M
gfzGWQbwR/YzVkqrVEUiKzYOGvKLFuCcCewiJlTNEtRu7MkQi6n1Dg0llkBhTlRcpIHi+f3VIAPQ
v68xpAyf845gFIJnxTdC07i4+2SczDtbgoeDnhXD7wQ5+FeKMsC7yPi1DHGIGOPrLEcHawK4aqCb
c39+p/+KiMjsxql+eqPOBsIYaNkdEzTi0nXecLIjP79U3Qyg2yfsrbo1Ukl2BUpdfq+OhQQpbVyc
zhCOozdBjRlbJIAjQ6BiVi1E0wooQFrjKPthpwuHnsEV16gfbyZfLoNb7nHlEd/Pii5AWwLSjw7o
V0896zdWAR1qdmkenq2+pK7KzGqaRaNAgIaO0veQsT9AKW1KzKuSOwrx7blpOSLMbK4+FTTSNGlL
n3k+6cKe5yuYpyuSP3hx4q45/dMNZRYlLQEzD1KGnzM7LzYHyanlKcr/MUd8Oy3Pi/UzKyqEg1x7
R0L9bX1XRhzwbR1Yd91rSLiUmqKEQWI8GWx8C4EVABCY4HvNa0APdH3ksKc5SFZTv/4iwfjNnSEq
PKuEKLcJWOCosipg4sqE8wUZFYcLPEaOUlNUTGsrp7N6rAX0auiL7wSx2EzM0BEI+uDd4xYThmxH
Rtd3x+jm87Qk7UcxZM0wqw8xbvIh5HUAQXV9Fx1UlxIJpp+eiN9yds0gjnPdmKZcqrEnDW0m7UHN
YWlP0q7aLX4NsFfj0a7pOFqJh0SOfEQiXFWlGCi/Us3JKnoVIXf8oQenJO8FglKRP9aNLfN2CHu1
c1mtyzPq5Ovx3TZXgLtKj5uZpBRzBxAzUnbG4W0MyupvKyZPTBkvBS5hCkw1y7dlsmBO2M1NGsjJ
+upkd4TVfu6RKrp0fWmgi67l75F3UpQ9anTqWBHZJaD5G0xXASOJ69/sT23JNzCN+1HIl6EEkMbu
QF/dvIPsrwEPjpVJHzOuiWK1sqIP1LY1homfyVskb0UBtQPD2r5a/JG016Ogj8EoXz18vGGktF17
j4O/grE2pbfANG6W58NLVjYklgdSQHh/AdSFO+VwcJazaKQbvB+5TspYfwjgWUfToV2AZJEmVm8I
O8i5BNPTkxrmlTvRkwTXgmpruHh5I5///STwKOSafgrw0hd5+cIdym17i1eodFd7gaqbVd/WWF16
x7MiVnVMlMAMoeKXe2u6Twi5/DckSJgaW6CoAg1gpl1Dt9Q1XqOs7lMJMwXkP2xYM4z6hN5AW0gn
dV9K0DEj2yVLLCJLioP303iMJ8cJ1zeLIK9hAV1H1E8UIf+Xq5DnmqcpJKn5v4RaQwC1P/z2Oqc7
v20oXTyqLS0ODuzGMaeADZnjmVwGdKMk1tbI63Fa7/eZeJrxyCY6ARm0ItrWvaMyPYCxOTN1z7HS
Qwj30VCdWNNkd6UqqRJM6IyrA/RfvbcpWGURnaCs6lMduvxr5QKVJ7BI10EIHH5TOrmZ5dVFIFWW
F5waPTu6AQBItralFN3dvoky7HgvRyN8oliHn8dhyd+jFfKvz6wbt9GwbpN83qzlOYybzMl8y20j
X4WpZLXBKTdkcvBeYBCk5XPDvu4BqV9MopHn8rHrvmpagKEhEjwIDDEjNOGC9XaSoKGgMHW2Lj8W
X7v/7DBhw4O3/C8ie2O4TSpJCAyRyuiWsX2DjL221dJrryXC7HDEcdJwKwUEInYuRyCIqe0rtqHF
Zd6KR2hDpXgvH/LjaBDT0Ai1qcAOhOji4JdgD70uLIvaiWDwSk2xc/5PUxVegOpaXw9BxftF5C44
8P76Asd8yuypkMWpL4Bq4zBbHg8uw7yUArW/IwDdcFU95xHOtBZOs03yhjldiw+Sr5v4WETTvmdh
MniDOspIU3AGI0ophY0QklBpxqfbfDFoUHLMjpXbj8n+G1i6cPak3VqoZ5XdinAYKN34bJp143aG
cU+ALsXQtosB2M1mB9Vog01D6uv/W7p4GKaAFs1UMAL6mLYqn19WD2iB7+8b8zQb7u8YVXEAEh93
92bD0hczBW/MwiNZJ28/HEjiR+J2C3rtOCYNpjc4Je58zwk1IVeVg8IvHpW6G6RMEkytR0UjInCx
g9HvS29B8ITYt19un4I+PAeoBFF2oD0wgb3Rj/rU21PMRYPIhtKdfpewCYuv4sREEVfgJoh3mdM/
3OsT1pytSELpH4vLAxWHvQZzZv3s/PtWYwMjhWBXDA7Eqd47h6gnqpWFV6ymwBbszEzrpzaMBdur
724X+2NLkWpitcqGuTtrjfXPbSmaLZju3ECUkzIKZvOQ/g1eEeAkxGO4JsGyewB1+wF7bgsRaYl2
xRm/LJPCnDVrXi9LVpLB3BqIDV3FUuq+Bvm/J2BtRqvFN9Gs4NobTkBwN1xmGwC3ddBfb4UxCwtX
hMc0SWtytS4fdxRRnZaUR/f2cqXZYNaGpPAYtTadnrDUm4rNkCW/K9nyqAYHNIDU/M+S9/gSzHv+
MdZsULQIBSlfh2H9TeMKY2bbSKKR3NqN0/32EsJYUwceMbGhTNCN/OZM0AGvQZk64GOLRNC5rKdj
6xq2jby1Jsh7yz2CZR62ZbOpPcpEgglK3mD0EGz4k/2rdfb1zaU/7bBLYW0aehku+0FW9aXWefCh
VRUahAxY5Owl2hlWLKf7C3a2poK2gCuq8OnG+emSznj0eA6bqgZKhx+a54SvDpu5zXjA5p0egj7k
njLE1PLGxcbhY+eh+DfqZMmgO8LlqToAbbY7nczuvEXpqa0sOfvFbJ/ax49YPwvsj+VwoLXlXGLq
870Jx5VKb/njDbQcLPEWG8VmOMUg2+LMdEFFRLyqdmeBuVVJ7MYXpKOMLSizizqYdJrtx2O6Fe3+
atJrPU0uCEvwvXouwpI2jTI+5Zs/7r6Tosx4/NtGLqtPSC/DbOLcOSPyJNaMrk7b3HRQizM7JWrw
5XhHgB/GlMs6Q7iQP1KmueY9WU7ODYvduEfcRiom9Mg/YrAmcrd2ptmO8wkIYxaFXYjAQ3l0QZHG
QPvMBAF733ChSzhfnW7eMGJtE+091QpdFBkeD2iSll2p7LRfjmG6Nsb+7sLxEXziUwjFYNx30+DT
4F/VQaszuwD35TffYSYvPx3IPBiI0PqjvEYvHw61rTJJW4bquKaD5WK+X2s7xA5fv8PPMwo74sFw
6R2BD9SfJNvrf9QRB7EGOtsN9L1ZOYDK8jPSnvIS5eo3L0bhSQ4X2G3qe3DpB144oRbghYO4YgVC
ml5TEOQu7pTPi6J5uQriQGdipDzDoaHf+2SHD/3VgRVKyDoD38bawe83Oz4cJ3JD17BZ3IS0suvW
2IrmvFSQi7RbIkB/DuVMO3P/WSFiJ9b8EvXfw8iZGohX+8iELnjx1gjyomfPOmgC0i21fp/tVism
l3X6Ccp8kG9d5Lpvdo8FQVYgXz5m+jhO5Rl5uUotTX6VDF/u0vtWcSfwLjoY1gRPKAPAF5WTWaRa
+CncLJvbk/k8gG7ptsqVXbPvFgudMDHgXCeVOt2g/31oHsaQhww/Yi5Y63WyCdRFrMA+yELGh7mC
/VURkLJ2MEyFbvatSyBm87SJ8usWJpkNzOgkQZvV0xySvPsqx3j7XfgDs9k5pTgcolIKzhg4+Vyy
lm/CmDqECEca5ehxmaVoSftGLy5hIs/tEZy/q7ESifLmAaauIwxlCEsOEdsFRBinU7vjlaPBY+hj
5I3M4LQW5QN45UQpj+RA3zBzK3MkLjBGAYmGlpab7ZbxmzWRsAq5YJJ2m5DNj71w35ZhSXDds5yJ
K9FQgyIKw+whaN1B+Q/+/JMcTuVUpLTMhD1aAOB3CAl6LNS4bf2dMuDmp+WLyvTVuFSqjAhceIHd
c77ZfFRNQq7IUtLJK46FE1Hisq3w73WTa6OK7NOdEtFUfxOferSN9q1xZaYrfWuVohy34VYiBGuW
v7rxtwCZQMP8y2ugR/yXbmuDmvfRHP61hhoXqr+rHUiU5YuUxinrjyF/nBp1LlIwOkHUopwjuaT8
N3hljVvrwYqRWY8hfSZlSTgGIj6cxC1Rh0bj7L+qprrD6n7aOADwsw8/CHyflt7udyjBOyrtErcR
FMyoCCJOEv1/6X+w1Xd2+pRnlkVYM9uSsHujUzu6qg7Ns8Ame34ZybmI77lSlwm/7LCbg9Z8uvzY
Awbp5x72hUvAi49jsV9PMoCJPrapgQEfBmPNOmB5Byn8kE1/h3PKs8JbPxspLT4rjoHda4OYIulE
fnF4dff+C0L7Up6JYsJ0zvcmo7c0vMRqmAQ6pwWe78he8xXyXMFWm/cPmbbq55wlKMLHZV9N0tat
G0KpodOjL0SnbgL12B933I2mB8hZrdh0BrB6PA9s4cM0SE6JNg2PpD9WGEibt1EUFsXNCk3D5ufa
xjVt7tBqGF/meedAR3rlcHiETPDjoI948LvBitETSnpaXpQy8KesvTKEejObFGqFN2hFTcW6Vkhy
IZ8SBDf57OSBx9dhzt4s9KrUtK4Oh8bW2B1sDgOzj0Bo0jOX6eLxDbh8boz6O0c3gDm0l4ASpj08
CMOJgp2OsXfRufPHg3u8dBosJMZw5wQjR5y8r6x4Y1jVkhv8X2XCVb16bV/q82yJ5kEOtA85Ox/c
B0lEeWrbEcrjHmKymCn46anXU3BMNIVdk6f4FMjWwtyDGLy3M912lHyLuKz2LUYSMG691Qez0K43
0B4qFIJ9LfnZcVHYN1Mk0DNgTPtG5FqwbNgEtG2Xoog8XBMrhLv2O6a4UQIikYtw0Z3h9B19zzZv
3kfj+TGnd7DOLoYxpUFDt9loFXFYuJ8XWiTvf/vff1+gEdw5meQ4BEcVykO8Y1lzRBWs7AXO6PJx
oWqImYQemxu9Eqm8+VFVWoAfgemRQ/HhkdTn82F3CfdeEo8tC1CvyzEUg7tJyv4AB9EKB7G/poT7
rl//lKkBL1GibVObtdA9qhaFCT9BpFFl1M6Ma/HhxjQFvT+fN8IpRH9cFirsZmbOI58ZGZG/LYU/
kdkq6QlWzTRvobnybtw5gp9fpeSACF+Dc0Smb97ic3hDDoWhKNHPIN8MIIc0lDbrufWWK4ZDHjGu
5NSFGbHwHx0K2muKM36wzDYP9hTyNMMfmqXKB3URFTLETqHeb7Cw5IoQ4T99nIC2K1n7E/PiHuxb
7ZV94rptjKA7BW/PTr82UUNpMP7wX356dp1EVQ+zUBMI3oB2l3v4xx4KnEtz8lIskNmWZQf9L5zG
IcT9vX9zB/qug2Fv/jTiKnToMUVA6oOJ8xsegle9LWeEkl6GMlc3nDm1qIxipuoy2jyG2GxZ0xLz
/7tMiHIphHXmt4q0bn1fztfErSQXMhSGCH1w311G9YiRh7K9OKqY3ie3NwV3s1Gv1DahXD9xGvg0
gP8yG7s77ex23MPK+nUCcjEF4KhB8lGxlmOWKABup4MO1Kw5UfoFcxHKaHFGJdNCRbNBrIBY8ukL
guAtFhBiUgXq6t11NpAgUuK6t9AXNl1CimAzNZSHRvxfx46MJWNEBzQYSzpioaGyYcPDLZn1MV81
sRvTkR45u8HFd0/+/y2z3U0kW/l2FHeVF98nT62ADrPTOJnZ69ETKcLA+iO8r/7P6WnVsiong487
GgIWsoWw1KcRi7sEAfWU9WEnCob1KTnrshC9YjTHVlYfOsbsf9CdWSDf+7O2nmGT1JCkE4kcR+D4
/oEzCDiDhAI5r5v7Sq03z0ToqKEsTuPgE0qlW/JjsIQdJ0mZyOoqkfMQl/eXgj6b92C2fsKd26Nw
QTsS/yoCRs1hoEztoA4YNeA0NwRk3rsFiVxNjCm39snyqxySYZdozusHyKx5G+eadlV3UB884Bfb
eWzFUdLpBUbpdYVwtGNuAdN6G+1V+D926Zk/5RBw9FH2LxwAut8wC3dfrikyLO/b6Zitcal2JVeV
ITJsPBHjLcAQYmV8WTcD80AwimiXspu2A5t2ishaVD0wmbfLZ6ltH5urV1Z01zWXthLAcOdVdTYI
QxUcS4bgy/L3yoqztY2PlWGyCBJChEsiT0jlj8G2rALMSPwcsFwcvTTrvxMn9EnLgjz1RczXv95K
CDCj5G2+Lr9xZY0ZYF+B24z4S+flFGrRx7cs9Xty0TFSxRNHCYB3TlKLBkZ48FO4N4DQHAJMqR5w
SIfPmFR7lOCjiuJnL+wWG1d+k0D++bzk6e9h7Y8g1HRFuwKiWdq3KDZrYSmCrLepOYyKd5+XhnMj
H+ftodkhxYI8LcomvohLv9DXaCl8s/o/wI4xm6cPphvGqN0Boz/oRrY7guGwm4yZQ+F4VblmtVUZ
mEQftQguu20yg79ffkocniyDMs6pvBxsWhZq8PmF9POKChkPki9tJtdPaExvHPUg4y7tf3cgxRB5
Sis2mruniTmZxYclEew/PHqi7skw2v8NEJFVZyBEDx38F3AxrH9qpUhFsLQeL2xVQm90ezSxiEFu
FXkMtfrv7kXvQw1x1S+5IxD0PKh3eBGXJ3WF72vHUmF1HZ44o6SX+681GeWqxYSQHMlqiAt249tL
tPzPrfrc9DFBD5oPDZQf4AEJoRmLOER7vGFsTu80UUa2Y13JRdMdG+bXGyra+3A03eNJif8629uC
EZ0n4QrVyd10bCRt7tdJaZZHPGc4+y02u9dcZrW27Ab1+ie/nGv3/FgE8ku0jhnCNckxeh4fSP3R
XQQEvB1bW/mPa8IZaCAdgF9+UCYfKkbc6njHls1woUV7J03BU1CerR0EwBQSiU5k9be4x/BlH5f4
zLvoj/uGgEY5O+76PODfsyQlu4SVv5qGOdUsDEMQn7W3YMcfZHSfFpGPPwJZOxdmK/6lAh445KxV
ed6bjdDiPubqKMx0xaaIRGKZlQExIPmRaXj8l961/AXVjHPHbcVQqc3UUIFbxBH4BJvwuOMBvcNk
Fihc7Us0sDvwVreIP7+jtQKx+QNK6sV3b1aHIyRYvXns3jH9mxFs32BSCk1dlaBSgG3nBOVQoAaD
uF3b6FVFA00TFYo6co6eLaY/Mj3RP08zeJnQgybM82Lj5gO+JgGaVEbAe+WS2uO/WGM5TCRxphqa
4rVS43cL26nP4mVh6oGROCVi3eWNRq7J/AWagJW0fPDHg3w9ofEvG1LVdwrprL6UQYxKjL4c2R0G
rcpMMPwb12MvT4LPRlwIWB74PLgHpejSUWyDG0HxAuCTmYEfkN0kpniDXopM5FB/Q67mHrx0DLQn
TUJ7dS6VLo9EvLSGu+ytccUJ0RDRI4iGW17vHZJ/KUXyNhzoRD1+0VBTVgM8eqySE8qtkuNsJuTN
nwcVjQXHNvANSsXN49g358B7lBuOKhOVNDq0oYDb2xTOnNWGc0qCOxqE/r6yOEYT/3J1m/EE+9o4
nG8/03TJZCFEYoZ8xdvs1/odCMj5UDiHmpAyX5ePOvmN0LJqP4TGmb+Pz1cBokqZ5Pmf3UHjOda9
4AKzpgfTnd+6iMmCoeiLrZQfaHqmzRNeVnSD4xttn1+Vzg+vVMv8wbWejZcWhzDrzhx33ViPwDR1
XmKX6rezpF/vxv556Rs4LaToCLLWDEAhylJP4SpBIOGEtxImwLZSPsvHbBYBFbwvLdvjuwlzSroD
50xXD6lbSCIaAVmQtnKLlGJwqs2LKcGZXkCIzKu4qHB5sIIt+EowcQvQOKnR7KJugoD1QzM6mb5t
n4hb2Q5n4kHFwmgi8IVXTNlcvjTZFuzLNNhR5g5rcbVxpKvw8L1hO+uI7I13Q4WeVbW2R92akL6t
8kq9yuePGyvXwZiBlm/YxeQ9tpi2DHzl8FHyCBeXiLNLyve2YqMSWsvk8145kGgo/K0LDfWqrJaP
eKnOjxaTN/xnj9j6VfjYOjT/7bFtRVuIdRRT5zo0d2sqO++gcuFEbjOknvig4TpBinP7lnPJurr9
AJEH+MsXRL4+R15t44wFgV2JjkTnw1x9WyETu0PYd+vcMhGl+tK4NtapfFg6u71CT/lBcr7zNECy
wkgv4MJwTGsr5syQPo+Tmx2U8bfktdAVpuZOvWvtH8PdYkc4/iSODN6xrG0lXGjX/VxJ9TwjOK5t
COJJ7ZGaB0JSazs2i20xfek7ndaOF8pqK6o7L+B1RmfAwVUR1QGfF4VfVY+r7VhWCOKqbts2VUg5
uoy+AUIL7FpO599M7wJtqyDds4i1y3kvTMDbY/yp9IGR73wbzD9G0EQ9kU8/3hEDwU+A97jVpHxw
VmetPO1/jyCPjwAc5TT9oPXYjHDfxaQyLTwIE+rxBgfwrxriTYS8ekr0FyU1hvwZS290Zdud1V5a
QDVKO/TVyP/0O0IJFEq8BVChUkpxVzKN7EHRrd/i9RXtW3dT+yy3svs6RoUlXniuv2xlC1a0vZcb
ZtO3o66brfeCOFKeiQ48h3SzwEer3lOTV+y6sO7707vA8acCynFn+4NLYY+9aRKcC8JoSNKjvreL
FUjW6QxSK8oY9n4AC4TxmyxC2qayZNUcjTJhLWsmY1PVtgUTuOYoywv8yt8ln+duade87BNQ6tgh
o3HcXPV7q+w9yxs4JMdbpc9nBjFOywboQo2zw+xAyL0dqQY9EZzUk/RoFfQdKywOHAGuCegcuUUu
RrmoKqFVxcjVENMfJhhGBpdtSqnThUjU1R2xjkztTmTXIWBovoBKE9gGNMnOTMYArvSVbJ4wR2jC
sQ827sVT1sSHpNEbXi9L+dgieFJVfwGgBUcYn04Ynl95D4dfxTxL6X4izNP6wIK86sQCF3PMEseV
M4NxUOfzskq0amofAw5Tc9GU6CXaKxRRIGn5AR2s54VC7T3JQ9Jo/0rRhnG9fCZqabE2bxcn5O5F
WXJzD3Hf08d+xmqDSnpATCT0X7Kcl/n3VQA3Tl+3o/z4b/Ce7qcVep+Ew5XOwqdfmDAr9kBujWga
AQHM6sHadrf6wljrh4PRZjuaIKYEiXETIF2tzpdRydRz57XAl4Gnx8YqMi6eiDyq62938XfTATxS
2F/oMCjVNf4I6huM2X/zqWSiNX1vLbTwSSvQvFoZA5FijJaQy2PexSRgfrN4utW1umFALDTpFD0A
tuJ8/mU4CVMVtaQLruD43fdCT0tviUvgKkHthBYoAT0tdZMZZLv/KPil/HIl07WYUUqIAg0oGvei
jQQw2a3QeiYaXzYUGZbHsn6s+XMxIhEhKvpiN44GiFZp1ONZKB9jRyA0EX8R/vms76jhgwSVYLtg
rzojg54ZaaWhmWnz9wUpvjIyM/ngfACG4Q4h3F7yPOqIx3Y5iIccfwB1wSQF2+56uLspoQa6QHr9
ytoyoq6AF+neQwQ3To/jSDTh+DqQzURPZpYpvZNjMN/OOCZK2nKlaqToPd7EflIbF9ksuHwkCj1E
+NWVPw9YtdqK/XezwOZ0pboDwJSlHniubHYJRD0TpMViCRN+Xp0M5SwLSk+0QhQBJEAx1VcUs7Ll
4IOKPnTFhckIvdkz0s1efMuoqmqdFZvBLNk26GVF+Htl/ywft3vb5FzXhguHsxOLXrZ2lfyH3pNX
Pmns0qPK1+JOjDL5enYMVGgiLFSTlzsqz1RfLO4JQzBvmtQ6m6yauTyxILIH+1UBLGoEtpSiribk
1Kr/Pgjx/crhKIkdxT+JkpDyAU9IGXDKxcn2qEliA+L+J7NGW40ntYEI6gJ59I3EWkcg/OqZmOkS
VfRXSdXT9jLe0iBI35SQ3FPLSi61YOjW5Th5ob08kxIZexww2V65B5i3M3LOGudTj8vW+m8JcSDW
mu8BY5MPvzoCVY/mUjBYXZdhW0ly8dnp8G/fPUnk2ksoBOdos2+qniXSU5pCMWlu65OG54ji+VBd
HrNT1iSpqFxDI7eZKpym4n3D4dkB352vz9caGObEFnxmzNWDraBsFG92kAOmik2WjPDJNFHP2UlT
I//pfG3HjeYrSES4IgxJoSou39hinQrelFCdY6+PhHd3tj1ouOcMbWEt884w0umz//qqOgwcZjyM
Id4b4JartoYQNfh7XPKm8zHAvfPEQgFWYMKgze/vNA/JlwbqVFiRFkpXvA+utEpDAWIvYN3n0beB
pgEQWJ43CLUOjQ5ssr5tHXkCQrOR/M2803Xb08Umes7HCXA8eUsk4HdVRQ9KHYMZGtMI2QRJY6YB
WfW31l/fPjMsBOimf9XDqh0t9trGaCWHyNP12IBGR3H10DLt+Lue2UwF1X7XBAjbZjTR/4t/91U/
43Yw3cjAJ+HNT/kHIxrNCyW3gXgT68QC8FZP4O20yKXtRcF2rBVokz26LnzmXrMtMaxQEvqZxyXC
/yqRKNi2vADoHbqXez2Fj3BJEUrRSkJ7KJqY6Hr1AYsfJYlfVL6TD3/hie2KBeHZYqVuBKexjy43
UrtayynuflOMG+IzJz9FE2SSiO+tQ5PQSsY/Vn/x5M83QByWF6u6hqWJ7aDE/W72o0EsugRAGb3R
axgC+uLTnqMXSZmN6kuyXcfAhwisS1u7VDcieXmEJBcMvKrIf9JPmoDq8fhQrxXPH1VQ8Wg/eZWQ
rM63GXT/xqzTzZ31SeBCXDFdjF47Fcf9roQJ9STjhNvjyvNylcpLe99MFXiXPCP00eyP3wgd0mBe
JBO4vD2L0YSnLUVWeO+yxGx1qbu7Jc/HmaGTKRso0N/ZlMCmVvcrLo4jS6ZSX9SsaGcIZIFAJiHo
U4A9EUGv3BnoqbUaCyvOxd/ZgGM5r4GUz9K+dv9WzR8GUY5ySR9L7as1PxgF6zzjyyb6oCjJX5v/
l8SooG/f/59uuIIrIEWmjse2SiP8vuRlJ1BaV/HHtN9nohLxHIWCagWp/CRQpFpPLdDYZJLaP8hZ
jQSHI+j6se1bZ8csQxIedpCd8E5RXUdf7r9N08Sswi3x2Oa38QSzKf8R00zndfK4/Gugz/eLOo3j
G0ekWDmoTa65SGsqGoM75Sj1nUww4jfXOReYkOORguROtjW1b0ZBTnFNlswVWOoYacZsLxPZlgWl
zfRHc8EA89SFN0k3Ytls1+6dZ4aMarWStZyVbwGSjXewqc4hi0huNlOsiqVGDZTn2LaRyRGaczb7
5og8VNMywwX0s3Q4a7H592vrT1DBmxCniN0k4aCyW2KcEpozQXZBvTO+OEurddcIALPTzNDwly1i
Xa0xeTTH98Uk6m8bu4rZEnUlk6UkfKo9Nff9YvbC1Ce9WsrPnxBdDbwxLYtOcp3PpFK08khOxIH7
VjJhEZGtwyPnepyAiLZmR46GOc3s+wF7tE1Lj6akj2uUnDTLAPV4infXii4D+RklQaRnnqswhyXJ
t96HTmhWbTKsCM6vTXpwVhhJxnIvVCw9p0aEr3FGzMdZ1roQJ5ZRgcm1+GpRnCJ3kqaZ1whSnvxa
rcK8CIAq9YyJ+yx+/V+mJ0KaHi01HQeCLP7r+h1fA2PsRkYlU1/0Zh9kNsaysh/SxsYLy52vxui0
Nz4gB41ROEsp+AAOSSBGhUuuOEyImMUj4wCPG32yOvp13Bt72f/ayaid7SmRxJsrGEN/I5yEa2kT
4BNKD6Yf+xHArZcHgz5bqgxtIyYYYK6A38BL4iCvII0vsHj3Vo9Dbn3omkox7ggIyH1JA6ocr7rx
Pi+QZcRkqMPm/tILv517apmw5p8A93SQ36rfGspzSrwBMmivZZPmQ5/EJQBSsUPHPyV7IziZdmh/
9DWsZfZEKI5nSNa9UWn/xGzEJOX2TKXuxb9Y/9XZgO3oJkni+7zVfMYRdU1NQAKyVP903ut1pWbj
g7VQJTKQCmWzFwoDeDWUbZBNNmYs1B1XoGEZpmwfW9gRWfYhkjQZsZ4g6DAj0NwZfeLvgzFwS/75
Czkb23o+CHCGP4S+THaUC0skQp7Yz4nB9wtwYcemNCC+/aiZVZ8P9nj8kDbBAZoXly3jcmisRUOi
q8WWjmKymlo9dOcwEeMf36hi/ejfn4J1TIkf/gr3Vz+FJ74jj31s91cz0Vn7j+pVmZwRhmXHqTs0
LKVwdU0eoHgVh9XjPilbMqDBGYzxNfl9dr29o8mQ3ye7GMLpsf+FhF0UUZWHIJOB6t+suS3rwS0B
N4D/rBaZLiVlIXUCDY5n4WTan6JsA+qQeFOxbzlsA1I7xmPrhO5ye+pHRFmpW+WWvKZ7z2Pm6STb
0/UUENbny3BJXtIVWAhVzMmjxuZQJDRzuUTYqPCJiNqTN5V5Mol0Xyb0hsO+cLG3WoH/97BxltMr
+N1imKQrh2Gt487Ge2YoY+6BjUIaJ38Fl+dS2QRm3FG3ytXKYdh9UDsUWup/RVnCCShXenpidUR9
WA9hPnS9OASJlB8DXm1QVe8eQFs1z8kvcC1raQ8GTp2ba9DSLyzdeSSFQnW2ct+AuGcuZcgLIvS4
Ifd13CqDCNHvtTBct9lV8VCgdJf9Bk22rtUgPE+KvcGeXYSb12D6TaDlgkP/+cRb8x0BaGGtz3m8
kkuCaobxOZBMtOq2ya470z2cba0c8zci/q3+XUKNEVCxqUp0HKr4FT2vW+3X9vTLOVeAzopoM+mU
wQy/Y2gvcuEKJXbIbL0gghCYZqQODQT8BAkRHYrSSHVA1TSdlHeIQKJAJd5NQdXDdcytNbFANJ1p
SmGtxrgHF0N9YMFmlq9b28hFzQpSe5Q8sR+FP4B8prCj8QOiBYzdMeRz+J67W0y6ThFslB32Yeo5
LqRMvjJCzKh1IFEgjLqqJ0r39P3qwiZmLBIrerqmaCF0oWfx7AHs0Ms+zOWgtuBIZpxWYfyEe0P0
nM1V6xt80aPyXzViVOqi90AUc5LqnxVmXMyR/+0rt/6qYUge2sK8Bl9XJ55dHJTsZuDcaAcMYhmz
GwYN17Y5QgA3NvJ+UdUF/0+cEGKbbSeEvD5N5b3bpQXVZUs8Q0l4XnBnCFZmSurcHfpyMHcSINdd
GQ4Kc3QCaDCrtxqTX+SAib9PbDyrZS3XBEe53A6MoKr2RfL8b+Bfx5OcwtjmR/CfuXa+zjUFZZuA
XNLx+prxH14LNFArkLDm6FZkL12CcN/lR7BZaUGVRA6Kdd+kuevR8ZcefbZ/llsYyjn2iQoWkmqT
d0RYzTqY07gAK1KQILjd69VlOMu1o5mgHk8NU6AghTFm14Q0ZNoA9JyFsaNhz4BKx3vKSS8txaS7
TKxCvQx2SROAPHE2d+GtnEIX3xtX7gTENxf9rrjrE6MYSeCvMMQt8ar9ubh+6iB6WCEehexLF309
Y1DXGtgFAMAkmSOJ1F5c5MnUhe5gdWzEEHnttQLpjb++dkygCU6U/0fBWDFJv1rD72iHpgVdCgMk
QRJbXWyUIDnRKaWg+4NZnlopi8fHP8AClMYdyPeUH34/qYHzDOQD/fBWDbUrMuxUA/yvWhWeBSq1
wPr1KUrZr3n7adrgj2/tkBsIjWe6NW3xkCIK+QtVfh/ZrZe97RTskoH2lG/fGXXg05te5nIf7Rjf
3oFno1Fb22CMX8FuH39zSPD4G+FOmi+jpjtHuzxtXGztLQvmerblXAyBDeGukoPV0d4V3vH+rcG6
ZI0G0TNzfCuxGAOsf0P5/CbOjwKUsPS2T8j6t58OMwSXP0mX1B7jY9E2YaFK8chics6P40QUoAB9
g70pGEwa7oVUS7YRpyoOrzTNOd9DaD1IdgTk92zdGTTSNuaHzOa9D93c5+d1tzuaheFgCCdwfAeS
8IltJmnWD6kCaenJTcwos9Q0yJ2/6JH0QokCv//sK0Hfiy1XGVspk93HsxHRxv3wKf9bGBb89XTi
PVFH+6YDdHmFSXaB96UU/0Z4jJXAf9dNSzBm20KgQRqU8C71sxYGWVoxysNG2u+7Yv59iTlWK5VK
/C/GW3cTve8j+XRA8I1VQx99b57pwGfbgIDvzDqkOQtRwP1b8DuNvQjR5/i7Y/NqF+3Rv8f6nqUl
Vmtdk9JeO+vghyA2dDWv12UP8XUWmNrS5hFeNWWsg6bHZAJtPGIlfxzQ4n8sBpbaDIabXT8UdDxJ
ILIVk1TqxZuqcOsv72ZDOd/SxLK87YC2q9A0eY1sjjf+zgBhRSS7ongM5OOKmIBxPqm/va111dsv
mwlmcmsPnocVSq2vBW9O4vSBtKDDzpulIXMfI/32s6PHi9W0vs1Wte2Os+oJbprprPoMHEjecMhJ
94hDTB/uH2FdysY3hHxb680KAE0VaHRFNYAZNRSHLrLeXbs8ZPESL8dIikOD4Y1C9Ro4ll7an7eZ
aONY68GVCPeHQFrsQiuIlMvTIqyTq1bPk9fjNNjnW9KN3BCy04BNVhQIvER6vErmQIPANmx4oEua
ualw9QoGdRbQ+uSPhQjIbLLn9/TkV8V176A2v6UZD7KmBaeNSyxUF4DGNsdzVmb0UwG2oSLf8ju+
u+tmHYs3utN5f2UP/ycRT5EVCBRnxZWLJNMrXK4tGzzO5fHTPTmmYV765R5FxK73nEKaBTzAN7Ou
EpiXDDPE9E/0j4J/h8tUs0yY5bs2O7X9Xev2KdK9aHinnVmi5lG+4/LMyge5inbQJjUmjI7kfmRs
w53WkyM0ytaFtw2Ag09EP4Pr6GOobgBMI22pxqnlJaRhbqQE9RBbcsmmlsTToDSbePVvTCQhUaiI
+pOYYX10JNv9B5rmPHqn/JwfOMHKJfAjpCB4SPTPwFA8KHJNoAw15flAQwN7YYOg8s/LUuucSi3N
dEuHPdpTrlGmUY4K+5R3Q+rX/v8uN3LDtOzUA5sr+HRzBMw82wxUm5dmtwXAA2daWILIpB8rUqfk
9f9EJu4AChmhz8fiw3L16Bcdw1KLZCsJhVpwP5LMCdA0mbHFeOWpLuq9PLSaMqutyWEvDh+YkFRS
Sulgj/mQQTlFxf2qJbJuDeKECerpIA3fjJMu5VXJicV6Fk1txvvCDTkWiRS2NXDQgWqdJRCG59bl
ObWzCGzsahkizDVIxu+L/TKSO57DMYpBwqsZ4Ur0Y7AJAY1nr9UqlJ2F5IDE408Fwfg/O4bs9ntl
TEw4Z/bxU/LCOAV5n03+QqkA+aZDMF0gbtx8Oaydil26VZwqIZIHKXXOIGCRksJW65mGGqf6Q6Mz
SnHzSfqTQkzp30zoOQ+LkHaKBEzshBtjWDCir82CI718IyhWpTdaVwLG0EcJsZ8gcny6YpQ02s7x
EYcewJ1WgNWKUwu/+xCha4xVDk8yNwDriYbCaKaDEWvzmoOz7T8gTIbFI8EOelVXaxJlHzVOCb7l
+42AZX/fF/7rM6oysqgYN4JzO2wG0hsl3He9lap39tvLWHFnSY5XMhfD9Je5ZuFkfLNeLziMk6T5
INfACttMC4CwSSmEDLjcbGi8Wyjl7Mhcs8mm4g9GvacUSRMpNMBq0kFYppvfUc872669X6z2ouO4
NwesVEYn7mn1XL8WuUewWCf/DFid3TTJcByG+b+J+YLTQX/JkvuKHSK4RgxaETmQbMyGnGvNATqW
/AD0veA90QViTOa9bAn47LKq/Ac5XpOeC8R78ct6cC6/vIZ+TtfmTOJvgcPQCxyD52TaDE5vvJsq
cOjK+dxMrgS4wojehzpsP8UYcNepvqM7mYTbj0Udgj1cs3Bcclq12CiZpTRzhry13U14ySRYb5uB
ehBTqtSs/3CLVROhYyC8putJN0ZkgUQYenqElDdALTLexdxPqwnFDdKUSMnWB3c5hyj9AeP/kv+M
Wl3liTcJDyX/xFSDWzd0h5yJ3f2UsVMD+BjTXHHj6UITE3JuaLesr5pqNJDP5jKqF72y3DdWTOH+
cuXnubD4Ijbb7Gx2w6kavoE9WvanEXWxqCDByg9RvjaCnPFcw3WKFBsTB5bQT5KRIlO1pCedhO8y
oooWtBhXGpobn5dT+JmAaNt6hyYsm3Ad0VnnMjbzYFufQfpE7S8f/wzsOuhXSVVAPi+uovFwjdta
G4OCfMpx1svMX04ZqhSXSRBwiaVstqTUvvOiva5BKwEf1ra5ebe3ltbIUDpzjKCsLa5+JifOuRS3
NOH8E8BBf1rW4anZE5UtLvYFVqtWsedl64w37ObOvZrL0P3CV9jx5x4fwngOKzdys4w6e1bQQ/K+
48qSt2WCC+eE0xGWOM/MGzwirfHLa+TBL2GUhOJ6uiOFTNJznMtBDNIqPYxtpqWK0l9AyKMk4tHC
8Sf6KVB75INEOee0njsJrK4aduHI9IBGviMHOPsT7bO+EeuGsF3tET+iE3fjeloVIPpzmOpfkya0
LyBj2OoYFIVm7pmp0uiZ+FeIrdH+KATGx3NnmyWLBnIB+tj3nocABl2dHszmzMTM6zXe28Io7L/g
PruTsaDa49KKmbwzvaElFYEFwWFhC4mWII1TLdLlCoQVWCMK6EN4StWBdfNDHfY1KtNcteKVP8Vr
xmpjkiWp76dsHJNMDqcCr3SqGkMvrN5RJzooU0WaZZkrTmT+3vq+641Y23lmvlYjJi519HnbBk2Y
9jSkrHuvEQoGHwGISfzOTDf9MgmkLZv/FvAsfNoaezGoCtODA1R1hLtgKJPFFsp0zKEwhYATSQDU
lXnLLEGusKht3bOLf6bmpmtiThDHMgaMiBZRAuLSr52IZXCgWs4OA8QF5Dgiu7FTx+xFZRYzDQVC
U4gvhRwCp6hwj2wShU6lpzxzoDclO6LgprEvW9HuhuccJJdnRtgv8+9sUctCCOzlvSVMuwjCQ4BT
I3zgPnV97hKOc6GCjIYyTQFePo34rmALrZpLWENguQ61FpLD8L5lUWObPRWlh9OV/x5LA0tbnzm+
JOp4d9NgEY81iP96CJzG4CqKDgHpFs62xaWvEDy4TDtjhzTqcgcGtXBgEViisfJVEwsAyvyBhFvW
4URCGlsgRSclBsaukAWA+3uC/ZioXK+5mNTlYTho1XPSAINlAJVzjow23Az61TuZjnTaDfHfQPin
GSp6Er/7LT1P2ALkJGfPiCfdZq2pE7dot4LVzATAg+qNMs/Zh9jfPgeYFsrcogNlXha5GNYBE4Yo
uZ3YNw5GBWGstA4v8NvB4omUdVNN58mmz4/S9tQMNlxIKulhFexkxFJGAmk5lPhhGKsCRp6wr2f1
C1uSn6XvNYPRapXpPjUfVotJKWo6hDLuvuVzUIEq40ZK2Zk4iRdjtZG3RSsH/ztiiG/cbVSeph7O
mDpzyIhs2veG6VFqOSDtvzGvVP+k2Kw6bdaaf75Ua2/ZZSd9WNq0ork+06mlD9kjOOWdl+P2c3Jh
4DDWuSzPpTHIT6cOywyFz1jcdasF1JaVzJ24GU4Z2c3WjJ1nKYBIzPeigwU1GY0zlJ0IF4LWi3yK
yUeaP/+u54iVMu6thOicqQtvSsQ1ExbelSaK4mpry1RlvASHAxTNrzXtlZj0x2goI8vHJ6aIAVH7
pIBUQ/37wAo5yCPQ7YuuJ5ximqPR3JJIOS9ho5lGxeamxTP3j4RERtnOIK3JxbBomQnTaVraiWTw
tKb1FTbv8Qy1s7EYObMr8KEkn5WijhQcqi/JY132YJxXQ3S/QD6SqWgUwOPznAhQHR1u6jHf/TeZ
YoAqY0ud80rDTyzmRcHtpUgji9DH1W0pKgwZLePVNTEZa5EGrzwnHKs/iqZAmz5vlHlZOO185Ken
j6+A7VsbCC6Jg3zW+a3crpm3CAsTkkdrFeG7njz4g3F+drFCmouOrlEiE0Yd6DD8oQRFgLy2xAMX
fYIZnTAYd+SS9HIVE7BtuwXOOlWk5elQb17tl/7BYi6zW2iS1aHBQOsFC6AVu43x89Wdwyqxj0HY
2ogyBf/P58q+nZsX+s2doqereBwiPDIUNGsMwwYe4UKwnRPJpBL/Qp+1STM2hVomURvBQuGwluQ4
HDe+bdQrqflvoKNERa9kBMsSNZCHOU6AJNdaP5NxDjvySHlLEtFO2qyMAmNVNPSut9UG1AcRgt0H
k9n44tBjyur3JVa9kNNQamR34cw+6NTX2jz7mZOXrc5gJiK2GxSGD4sBIzkK1TO2dT6+sdM0ySQn
qX6JpV105mUNaEvFgBQhSa1TeqZueQJoOyVDp5QrBYG+t4biAW0ZQNiXDgR0xHMRR5f7l12/5pfQ
WN5aMMVDbnm2W4tIDKmTkq/XTt/4BYn1Oa4kMpiqSZ8IFISFajLWecGfeHqpC/qI1PyZLM67SLoV
PfIdwBCZhZMAWmUahOd76aZQHCjnz7RnhdNiScUp9Vac1C7SEMLRy5xd/uLCUgNhfS++5j0QAi1h
QMqwdqBNrKLlCuCg79ujaF5K1Ft3JOHGu4ym9Hu+1FtmA5Y/9j6yFfFife55ybe77xzEsQJR3bIc
oMOVyQbjfmOr8if+2CGk3uuxQd3v+S1/yO/KJAfAkuJPpI4FY0p1Z3KYTlPHOseKGk6SGwVeOD4g
kpW+UCGAxfhv3TBTvs9sSR6oj8ZYgJ2pQWcML5edXrw0q1x1JBSYNp+vKtDPZ6NuQ6eIUyA1fOA+
DnMUFOYyBx5zBnIVRshWxS2dl8DhLlUPF7v9crbOInguYqwo1/An96iQhSWAioJJWo0VDQ2ZQ/a5
MPp+txWlajuVLLGm4E0wQaTLX2ZOfZhSljkdutPty8DiNRdR9f2NgTVEWtL+yoNN7XT2Bdjpn88f
28ssENvcEbsQZQS1KveUq7BOz6rTaTEr5erd/Yxv02N5wveLRF8qS5cyMj34e7+9RqlhfxhWIIiP
aanbpjYX8sVCfuBxd/Vul0D0BQVr1ZtMp6V/Y7kEVG3jg+HY9o0KuRZXvo6GD0Qq0lY5htwbzYNm
O/PlATw0Frg7gWucAwQB7Yf08/OLIfornFezqEvFDG67fUpVbovbYL+cQ78Q94NIKMIVp7wihjz8
3EHtrJOpzhwnvHOqn3XsXH4e5IBkR/CQg5TGkk8dGL94CM1E96ItNtNnvleQN1Xx2fm4AfNjT54n
eOB5kFdwFz1iwgk8mrVCfa9h5KKjbJ9Z/Uh543dt6U9x8iHpYQ3Y++PoG0TVCSqBM8p1zoxnYNmA
KY8higJ4JE5BjwRWcTGDamNXCQdA5sk0R4EEX28KlJDxyeakgZpGjekcUUoTmiCzS4NMHVGWVHiV
MKR9WNWyLoGuyP4/9Cnr1+0fVqCULU50y9bmKOdjDD3IAiRSUgqkWuHxs2x0AQdfIMcdPwcwauZe
i57fdIFUC1y0xU4WdwVpG9Q4L/oEOm9xYOJ1Mx9OKs0Df1pHfNnx0DjASFodDVuzblymc5JLiTx4
udYa62WI7oW+2NNz2qGGH4noAqM0sNAEW1zdJvDlelvDaohr8Hb6eHzzB3A4qsiv5CkOBY7qo4QG
KULLIz6UEWsf/XovQmrZ974ndn9tGoffyovXc1ngW8GzeldG1t/I2aVuuhaUxF5UACbvdZcWKIX9
dyt9wrkY/I5ud406qQSPrea6I/cXMNld6vp+SitPk0bZhnLHt9jBQ5zog81bQ/0hdcTZeA14fLyz
cFqc5LRfvpuGMKTQXS8G8ACrNTLBNqlxR83vj6p8KOSVBOq9kqAHRcsY3k9Np3VBbVNGEfttnODX
kT8wtqRbMHw6ykK9X4pnmlxSfjQvn1uPYorAn0OFaRsi4R1ALnwhaWGSBFwicbIyVLAYTBQSaw0W
1eXjqmZ4z0CavPQTRL16dW0UKbhxMmfArkWBsdzi7g0FiVnw77jMjIfv9yxmPm5Eleh+dpULYxgz
LTryaUCj2/axeGI0K5nvwM4p2kqEtxKPb6olDSNX+Gckj0+Pi1hcCeIEILNclVdelFJ56mTomLWB
ioNjKGDBQMdXLsyboJLlKZKbWKcBc/5vyO/gVnErw5e28RDEpb5ic6eRxn4siPEd7u7S2haE9fHt
HzQ79/uphdYf2xMgUMqRO3Z870LUX9tqb5mzgFDNYV5lowkaz5w8sCFOuaJpQZpOi5gIoKcwz7d3
A8NrKfb76Ii0ucXxzEXhwxHlHg5ybTEt4LtrafeYCkA8s247WmAWU1Ff2CeKBquGD2l5czlUcaMk
82sMjNsXKj9y15GjV+adgsJrasKlmXKZ7Kxzbe3OR8ZQOnhUjlC0jnW8T61VUL0mRZSaZ3cS9xeE
ay7AE30aCnZ1oRBpGQ7LkHybxwJbaSlh7TqSyRrO/UCahNTZj8FHlciAABTbCaGHQtUb8GpDszwl
3av/oZc+/inOuuEOrS31dUw3vCAzg/8eijF6Bs3vpKlBYfA7KMht+DaLuVpAOKXne6MwzMdTmsTw
PhbGQzKMZqmjLrT+PxDd8tefeFOmrVqImswQwa8PnoJuFWkyJq2IIaCLCaRCsnVJ3WOwB6oiJE/p
7JMyXZ7jeBsqLTeCT1fYdSJJNB6gzP2ZJIUTadudZZWmSRkBt6vXUUMNMvXOmTBxPgrINxQm/vlS
4DgRZpvQ4tmk8dVf6XqW7XSkCy0TibgBDDKZwCyRRo7j7lFti5vj6E+5XyuemUA6X6Z/R7iZfN3U
pddQiE+Yi+/jvUfxb8yniJ05Ww/8UU77hBtw5jTHLuHcRJFA5JVQiM7D3VbUB+jzuBSAzPq+rnwa
f9C68Bz9xpar8XGzhSDk0dcWhyA2YtKf4aawlP4WPF0whWEbCpEozVtKKXRQmy482Mp9WgfkPRGo
ZF+5CItoXuhmzYpYKFozhzNF5J3I+jm7dFj5QzEgva33d+R7/Yvp8p4IJa3WVh5Yx6dubbfpBbcm
lPQ9pZgGcLm+bbluMYXDNoCnLt26PNyBln6yP24nE2YwLu+SFQHTkueaRgUUgzOiIP+4mnE8V4DJ
1atgV8xoc2iCp9GzVIzavBFoRrrvCqTm12c7TF7N0HJvK3t2xSqCnrZhZy8K5flgKgCwAosfx+yu
8ScaaS351H3ibQ8K87JagHrzLsmjQ6ebKAeFBkUbQbEpKIPMwYN5gXq2HaFQPpSddhUe5esm5mLm
tOPPdNo8adP4LRsxOaMt6xCgYjU4nZz7MFxsB+jRLFKdX3VvzEFs7BV+lprljGCakej+g6DD6jaN
lmsdir5i3bvBo3QNVoTumetSnFYHlSDU6eENb5YnCWSGUjX4FX/CpJcNvu7lXIJidGp4HKK5Hfm+
U4LbcYgLVtSJ1HFQWQYOKZMUXJmZZ1cqMQxchVKah58oJl2A0GE1pyMnewCmGe83rnzF+rVO5F/w
xapMU/qNZxRni6Ht0QQHaTcC4NYKFW4vZOEfx6Nw2wp4RHoE0D2SnlcPnIhIgQs9YUNUdsBqocFE
jq9U2Ck6HCzAs2dued+57i3E7/Nxcuq6YGTHapBExw77s+LKwcdS0yBak1UYrbaLy3uxjnOt6IYo
8x6ChMQ9ZwHiDUjJbJzd77cIGkLa3YEPolc9Q8D+1fOy8ye0FPX4Q50DEjUhbCREr270AepgIWSD
gAKLY7pcSscHFqBPIXZPhcTQnBgNtCQogKmL7WonVH2G3CidGOvdLPfurkEh3PBbpjMKi2M8lnPp
l11f57j8KCFpfo3Tt1LAJz4UTcH7xqg0nkIjUdEvJGQCY7dn2Mr/brkE/NABCf5TbMsTVGJ/Haun
uSITLtyo8jEvxxH7ngIuFh7jp/38h9+D5T4aWiVhJkdN2+E8a5HA+kJQFbWe9k1W+q7h6nEjujTZ
KBs/f1K8oOCwjB5ZLleii6/OH+DV7rDan0qwtDytvniIFMWZKv9g3vK4mAfFclBbXgpIX8dwXTa4
MgETHTmMTDpt9whRTQ0DjFNgF4sG8A3Y6MM6f+NtFzFqt0HRwefh6rsdHyQTZzWfkF5us+FAkQ8T
87MwjEMwQRGh/F14tkzZlcWG6/w4P2+VWTi1nyftjcLnhSmaCEs0Inf7otVGzS5TFwkRqA6OcAKI
btY93mI0uj8lkHprNAiqBCjIy4jO4L6eVy53K0NiK+DvOTHhMTOuh5KyzzKvWimzwAWM/Dzb10Gn
XbkjQ4p7dgvT4AJ1rrQpHVb9mLHDxrZyVOdkJeJuQvzilz/0glfWncw0F9dq0ozxGfQ5llRa/LF1
HrfXSe2kPYgEm3Y7vhhX36j7entAo8FmwW8zYa0qok8LQyNGtiO79/z4p31nlfn86jC/8+YBSkol
yzag1iUGoktjAyajxQ4POIzEU4XCLSC5dq5meaf6nffy4CV31pbR5SGT0PZUDi/D3SEJyYyI2wXk
fvScAtCIkMmi6sjMfOfGdudT0J+7pGv43t/DbsPSSCU9dh6WwxVHgKR42wrSJ7U0sBN1uLBWhF7l
Wr0oV1tNE4rbXx/jwKi5xfdFotuQBy4uR/rbQJm6cVZT2d4hHdI3jVJMsLLBZwMIYIYSx9Ej6FPi
a7IssC6sQcKuXmdJ+yoTRwrzrItVDvwVGF2Ubx8Qw0fzpnU3u/SgFoVTx720h0EP/tjN+HMGTWYx
rivZfLJtks/PgaH1OxxOt6pHzOaXa1lSGsgQTbjy62Cm4dJoO41yyWKE15mnHZ8g0444ssKIhviX
KeuBrN+JLPgWPaFPyzX4KHpDfJ6cfsb3m/2RLbtS5bxfs1u11mEjqhP+tOlNjosJ5tpzpazk2hJE
8E0oM2gHLtkfpzpjRdN6fj+NgtDQqBo3UA14XVlD15GZDYcNvht+6oehq2zYS1g1xKavwCQrYSN7
Ymc/98RyuEEms3GgpWa3YGYULSk0EVHZaw9rEF860apXJaJu+MDF3oJES8Dluq6WIsV0MHnsMkxs
pyiiGdy52tJRWjhrKGJ4bfrtYfGZF/mb/mSAuYiuMrZrhAaCPjAaoLHjFOyNyhEsGS0sG/ywYmwX
nbc/Z8t7mXOYnWFYIWWUaqbznouICquXP2GkxqPyt4ICJavF19cEIAqkK6j3HrFr5uAkSkEijbsG
HjoGMCrm0nfNJCeSp7qWAgQGrZykyk7UgsIWGbGmtiWwhTkVIpxFVAk2DyalyVZs8s8X2jKhR7iu
7+4Pj56k6Ib4TZEOgxjyxRunUuYwFcliTBT3woYQ8ER2G0kQgoW7WCItQvmVOMHdqbhnqOb6hpH9
uM5dZxgoLy5MEiGeDwSavGvpk9m26IvaG0eIaqpVXVAq6sWL8eHzD19zK5l017ey27xBLoEcbj+L
v3lcjo2oOlw9eWv8M0d1lRxibIxYdf8dO9yW8WQcSVe4JS62soFUelw1iRgWuy1blNSbfCukac+X
NmCS0oIA8z4GJNki3bQJnd5a87bYxdRBWpGW7HkQ4e8YqvFDwccLRLynRR1w44r0Uf9jWZBcfTZ5
FMZgH2eCU4oBblDxNiEjZeBAUr2uAl0zCXsTtM6KGluXGfwbUgmhR8wlRiXoPGShB+NyGGvGlksl
QyX/2XZPnPkP/5TBkcptBUH5ACg3LmRt6oRs7Vr4repLtQXqyOimOUMCy4xDI0oc5bJ66c68DnGv
Zwxp4kUH/I9mfKvkK51Vav5roKquN7L//hAAE/OORZcPpbIhY6POIK9O2NREUuVcCfPr6xZIC/74
UVP36sbilNEskTFhEsL1JwLERtfQZ67reSnboiPsbcWxRqA5RJ6Y+/Lpe9gKt9kZSNsCwNV2ypH5
wCj2lhPmg7etnxiSl1VJBnhXZf3SI5swpWxhjM2+6ZHRqsSZZaoVe+pIsNmuMKQYxBuZ5TPdHK5V
VnGFsm1repAL7yd81Cxf4PBco/M3bmtv91a1yIQTp/vjMCzTlpjnaB424niIlGdzgYbCKPLc4+Qv
td1HnTZ3QZJAa2PGOGYQOhnXh1NkvKZV8RwyI+7OJcH6aySvwStz056sZGvUall77/zxDn95JrY0
+Ue8nmN563VRy5s/rhB+4FfaY2isaIlEOSAMvXcA6xcX1xi0vY0Dm3Bs4I4PSuGaeftgIYJO8XrI
ATs1lzOKht4mHptc3G5dOXUoQ43i27jKDZWTSzmjfBbofVlPkA/qzCFQV9KE8KFj+YstneOtD5CW
u8Y2wHn3sHD7Vgy3vBF4TdzUegQ4XZJ8WwlKZIqwmeen+RyzhQo3/B9gpNQtXgIfECln4gyd6YKz
8i79j8A4pA0kOMtA0oo8v+q7KIJpO0IsXi0WewUiCSP9bFsZUfQWVY3sGbEHo8umgJ0dMI3qQ6Ns
5GVTUamNL/u9LmOr4Juhr5iwXoGGQzbNFJSHvt649ckivVlg0T2IOccV2jYOqCvZBPqPtT1OFGfc
uI2S9FgtHG9s3NqOkawCAWwBlc/RLWOvdqt+ne09E0CJvF10zGZBAw20iLw61rhmY0l+IPsjBQm4
vKexxBxpHfa/GbV9v/YgIArruZoD9SYIg+0oDHtc/4LztGBJSPDy66Ib8bGUY7rpS7ktIEDy6uNz
ZrgcFr5LfKlwe4m42YhGPuGhem3M2hj96qiaTxPbqWlkNILgFwMt2NZlwX25cxLx6t5wGYudBaEx
Qh4OwNukcYvdOEr6jBbthSoN0NJIx/HS8fqi9iEDGRHEAIjauivOd6CKSZiPy1UcNeGO0jfrCtCY
6gtCtp2SLf88kddGiuUGDMW2cszXhj1mt69uZKpXJF6v51GitbNRJHvJf3wnPSHgZU17Hz+VTSjG
tYI7PY0FiNBrAwsdmKeN0ZDpeK6HhHRG36hOX6bKj0Zm85ssbVZN97U90cg1+ksGIViFBUXj0h5I
5Gny7i2+cjBd8nJZrVgkiprWjLKLhzgQgFKYvlrZ5nCiWTweSmu4lMoybytXsPuPWLztJbXrY6St
TJIK2Ebyh/tqs/plMFPFgZ7M6cMA0WddTUYqfEjynyFv8y3EKSHvgP67lajON96xW17NnydBvtsP
ngiO/tvseWFdwnZJKw/izmAjW0ySzI1jyCAZToFh2R9ka2WTjyjWQNNtECsFmwFZFXHXvjf2vxcF
KXys/zLnjrvW5lzj63O610+O1sA4+JX1857hNWVI2FO0rmS99FpycSrLhreSGJ0HbVaSqCjfTbUu
l5GEAAUW5RwzIY3wWb5TWkSBRWShQlfaUD0tpRY0h/rfs+SjBPv7zjyxthYl4VpAHlwPS9EPlki7
lw/k40vop0CCs4Sgaqw9GudXMWCnsMfVBQszQdmynWxuE+XBiKLZgmQhzpg7xO6/zu2y8/2vTadg
k/aLH7kzKXRWe7jItNSqbvvlKu4PNokGub8Nq8QyxcMsqo+IbRV65PYf9Dr6BlCebYfNGYEwNjb7
Oz6hreJwnqX2G5lpmQ69i1madJXiIpcrR+UZdD0tvFX0TKyHyvMpONvRuDqmpE9PGHFOluwmlL75
W35UTnbQ5/IEsHnOHKglXAPRKKRCDDNiRiVfks1VohxLWsznxYL3SuoX/BCpkBtcid56DgJJUPMJ
mUOZpUSKVd0h24roU29Huc48qad0CdNcrMSOifdglshUhYpfWRq6i8YG385gZDw12Pci7ycvDe9/
7oQxFkoE9HcxfCN/3lSlVxpw65nixjRshr6T3Asfk2IzyVT5vLG8heeU2HI9uakO3fzbtd3ETNz0
DR9zpRtQA4cXjwRKkBJS6xj/+BX2MJ6Nm6z6UMAwYTU6SxLmqAr2butHIVuZBLfFYbvlELA/ySgF
ujtuUhrTE2hhHzC8NYX0O7M2cM2yu/V6ORC7n+PeoPd3QjoJA2SD/ZgsT+pC+UoZ69XRcfF6Uft6
gz/ycB1BJul4X48Ri+y22rsaEY8kjfrcZh9JW7EFwKuGgwU9+Z6gExfGJEqzgwzB4ntiRuvlhfbt
XJKVn91Q/SaWcwxDyx+jgUrFDdaN0B37Yoa8IEmxkx8i364bECKgOBdlubNHgRWkPy5IvIyg/gAZ
TkrPiYjPOS9fkO6tpr+0cxRw2/TI+ZZ8Nmi2pfZXz6IzdhUyw72ZJYD3CTdCqJJsYnR0XDzbNdts
41j7MTfHNsthINs/qMQ84GhQb+2whteDUVpf8IkNZ3R4OYofOd4uRJsmsyCCtb5JFP58yiQkIL9n
33svwvgfGXSuVI1n2tnY5C9AiHZngsgXUVcaXOoIUaJbHzHyIk/UMt64wKaU9ppl9x09VIOXiJOA
HIx0Kjr/9rtdyaCkT3/hiB7MYt+eGMmxoTy0sY29eGmORO5clVl7Q4fcidhOSZ6BG0lxZRYk5tHl
SmMrrY7O27Y+gKPoGG5WwucVHNhgZ3VikWK4l/0gfhJ7Pc7mO6EJz0XlcpVTphcPnYVv+AWDIvMH
qYewb511AfN4JzKfYxofuiqR/iRbpFgi5bh9+l0SgoFbqR/XpCk9k9gEK+Pgbk/hCo/gFHaYZ08J
51TxlmnxvecoRZhctLWv1Z91bLJZD5cPaRzy2nHVx7588pg4b+FAyFm9OpTRitiorN5tggMg/PCu
kERXGEndUeGGMjN9L3nLai6AT5WnaaGSeckmjSczukZgXCULfPHxnEps4Vgaa+f6dAVgTyDzH3sy
3wAot+dr23euArqMa9G+W+VnjLAsp9J1AVy3sAdjEo6ePH/kZENzny5WJsbyatgNusozQseXuchc
ooolS4xDQMxLW08uyGg3ytHhkVKpbXBC+Aj0ht8SDu0zULWa6dIXge4fQNxaRVRwXyThqfDkyPwl
dL3MWbpeSv0kEebDhl1J4L59PY8HJr/27EpDx/ihBOOTKWCRdamNwW8DU2Ln2mn0LvGhnJvH+6cx
OpJCgaAjEYL1yAY9cTfiM7yDz3HgNRu9BUnKfbDBfW63RMShikwgraVNgIXKbhPKA1XH6mj2u8Ha
hjCZBQH1jcUZf9/dnRuhmgjr7Z283OD7Mf8aogRI2vczHK6zcQyxgVL5CWTmbPWfXqSq311shVSi
Od+MTCOgohCQaeH3B7AfQBeqPR5PuFIgsCEQW8OcnK5/Y7ue0eQcf97u+IjCLlLiqV4zMDJ2tki7
Xpq31+7bD17+MT0fuL6qT/tj/B56eWaqws8JD8Go0MpQmUQFZgPWm350hGeJrIQuwi6xogDZ2om/
LzAMNkPtMeZfmCnXEwst38VmuLEBa++GlurzoROvlDOCGK257oGDb3qZDQievRmlThgIRSahapdU
Af6iSyuvyXevjD3w6NfKJJkIhpWHuc5jd1F4exkVCMYar1lCLxRtKs1csKBsy6+OXkHuKEfBWitz
s9iAWN4gphvwTLyehZgJ98m1n8gRiLDe5wfPsDziYH19eri433R9mFrmV2cjtUVXLDk0qCup+Z6I
AVtn0+Eql+18+w37FQ93TYBjnYPrBrWORePIEodzB5EEaHI9pjfmY3L6OLnqe3aD+EzK451zDqsI
Xob5N0NCeHJKK5F4DOvCWOXM4TiQUJCx91hRA1CHM5i5UwuL2r08PI4UpzJDG/WkbXx6L0XTQuSY
w3HXs/1jJIeXqK3fniuG/AhIsIPs579PPj7ilc2rDIcCACsqRpkR1PMTJMQ9Yc4hi/4EkdQQnNhB
QqjK4OPNdJLOB04YmpN473ThCooIfHilvIztya5c8fABrjVyf/wxS1rmxQgDjOFnN8+wHf2ynuV4
R46JeECBqGHkpO5aHlajX6c0fOgF0Xu6CWViB4TjDGxXUc9eS4OmSBJAw7gbNdYsk6MBeQSoRtO+
QcBv8HyDUE3B8Iq5rTJtLL8CR1Z681t/NSkVPIy4yKn7nf9uYkhL5CDvO/TZ9e5XLRmjLlAYbjRc
klY8JHuS8c/JP+XBKxr+U5Khnm0VJ++A31zMVrxm3NTmGl9Nl0Vll4JmeO4UwQZv5CEsa+4LRjea
QX1akZ2VP4xZwwGiMjtg6IXnhe3L+OL5tR3+h5NoDrICpOCnyTwbxbgE0tzZxSsOkmGgtN8mstcw
Duet6+aqSeByMKfbP8pq20WDzjDxu7PSP9UHzIgOCuWED8Sp/AhGilQixn/Zj8U9PwHtVYECeZQt
lnU/950qOCzlSfKDknm/dLoV60rQ2ELOW7XN6G46dRByx3ZDZXR6HZxRqPhn0I63qWYyk6zKF/Ac
e+pgqjR+UozPYbfbY5aUFilajBW+WaCd7v/oQAYNHYICAoofdrfv7VXxDB0SAh1dtyebg1OUy3yt
1T8hcRIWxBbniVcPR8dzj5geRpha+HGvZXKFfOZEIzCJt+tBp6zb0txYUpHKo9cUDG4X1iYnUt+P
F2QQIwIKAl1neN1bjHK/iFIh385NbeEta2TQDorGJ6apXX4WI86P66JxPY9VpHm7+BGzJVwzTKnL
7Kaz2UJhiz6Ta+rkHMte2KZfcRFPqKCLZJ8LfokZETHVV6MQI5F9QUeo/6fZOP9HBewQ4BN3lB+I
Ud8Tz7IZi8LU/c89pWowCjtVVWR3Bq0EzCqnCPcrbEH3GZmQK6YZS57H8ieReWEFyhfyydKbXY9d
1siir+L1zH2r35xEZovlf9uA9BGvkm7MlveLpv1Kif3Jhq7dLos0CgCYGUhYlVqV8tkZs0HbZ6kz
xCFIEuIVCQIYu2cKG0isYQC51ZGuY/8KaRr8K9w83jNC41BEqr3ryooDl5RdEjNW/Tw4ZFR0ge9S
M6KC0QGV26/vvGHZ+TWv+reyNfHVh3oX/pZILf2mn2y8xqxMvkXP7VbUbNnkiOs6X8ylScpyg0AC
14DwMws/+DLsqHRTbZf9tA5pKbdgk5sTNbB2Zu2FHoFh21VspVoCKzBXeZ1aoFtuomZIEec1TChu
t6LHm6LqziEHxWIc+NuU+NSeDEd3x2TgMBmmdB+oGbqj63z2w1Br2njFwUyaQPZIylrTsB2PlllS
wchLDf7YX0N6dSDhuKKQ/4xHaADZL49P8Vp6lBE5PyR0nmePfpHc/2YCBFNSaVsXVssM+OrRMMHa
pnVRu1Mqu2kQBCFO9nNhl6Wvnr2HaQyyt82tjjS+nF1kT4jBXfAE03moxlGSSnmBSIeo6TIecHj9
EAbfQe/B8PyvZX1W2+IpzdEaw39a5P+VB7vqZOkSxl6g+HEYffsIiDxiAMA8xKiRVlABl6NA+ezL
WB/r5408kxd9f+j0KvTFduqxHTMzb4N0/ODJbbBxsLGr5zjxCooGyJyzvYRTolgo7VNvIFVYylno
7knT4LOEm1dOVa+CfSfd0a3Y0iP9HLb/NzGoMmJecp7d6Db0CMCxT0A9KdplJMXUaZqs7hUwh8p9
UmKFiec4djRivr2NYnA6uZbU2qPh+3X/LelUbWOgMyCp95qBfxxzG9xcuwMrA6P3L/8qBEf8gQz0
R8RaSED0I34lS/Es2lZJU76MYHVvaY1teqHNIC4lZ5Lh3JijpSEODnbnN1cD2Dw2m7SxLw2J2fM2
z9SX8XFE9luXdjoOkMOLfU/lw6YSJkqNfBzw/3UgH5efA0WFgKdLELm4Wc/l+MxWScnmNIgjbjyJ
FuKYjR3ziLIuSVPsHUV1t9ESPYKy5mijbgIUYDuLbCoeobwiBUJEiwDrnWEI+/iHWF6yJc6ClIy+
Qwb/ggpm6Y9sGDTq4dIicrR+U2vMcufPsIsovFLDgU0AIbQ75rXkBXhIsjS0lm6qn6xAIBidwDlo
nYGUYFMgw1HJzy3mzyYueSdGhrPkt2p7PgbxZeLD0ioOISH4HidhxtQ6ssW01eqHHbjtAG56iVwL
sfCOkVx1tml5JJDv2e+lvPP9SxLkFAnujIFd6hVznVsuikFmc+M+KrnRSJqwUpL1sofheV2fwYxw
ZbPrpla8zUoTimAdBpAuNKp9DJjv4UsxobWxI6lXQuEt56mO/IB+Sh/8mMR+jjB9t/kMfhkX3dW6
oUil8Gz5U9r88zOqydeavV9r/2Qv+H0NJqFUsMuCEKgm6roTD93IyE9dvZRgqWKamRoHcA/vXTLI
LKdYaRPFJS3+l3xZ9J+vWEiFq6y5y0Zrr/Z6O/97SNEzIwD9XqSh3c444iTsiY5tSBoFq5bOHFOA
kiwbsoFqyDGmgn7qFd7vx9Ac61OsdyRYAvEgRVNwt6ADVuLs8dUHiMoofbQbaIEmkgElwoD+ZD7K
WDXupL8JH7T3YE+VDOE5qiO7ndltUu6CE6w5gjiGevoUzNzcuY7EchFcPoGsFqXEiyVHOGcA0tej
44reW3ImffaKw6F4BaN//zmcS3puyACNuwPtFs6yXqDK5fs4Eb7RvdZVzR/SYEawohWCPqsUgFlz
nu6Y7pAEnSPFtryENqAWDfLyKpoYdYjyKOPlcytTTVSlAj6Kf1wVxIQbXJDI+CBkLaId6dKHiUbQ
2CE7lMxZXPcbJWPs+61FTvxwVwDnkavY4X4lGqMLuFBOo8ds5SPBuEhAIszrGD2b+BGgXyMVZBQZ
HiXBlzi7ny/72xhGawfs6UigqOIJiF4lqdbD/SoPAXx69UsxciIr2mpMUpKJ5DAKlsnNUSXO2FAc
aAY4RfcE2zrdIhKEREHj8NK4f65NW3w0lICCp2hyBKMsw3veli9zUPsWKiW3GBEVHFuFVvy3ifHn
U8SWqYDIixQRo5SM0fetNthJwFmgwhu49xDdVJCzaVSRhtYoIxIBvYNdIbwYsvRb9Zb8DCFzzolo
tJWPwy1jFPg3XMcARiw6r3WxhN/g9Xdbjgec8Y5gpujdGXc4ocYSRM+8v9J+mMduL708ajaiztB4
xT+oqHiWW6eREXJB2MW5cuk6+iHg05W3TMqhQjFYqVn+xdcE4Kz1sKMNkpLhTAl5v7Ocy9BfXmUe
nRRMzRBHMxFN7QhDErmit+GdSqctTf+JskIUlvhYOyqEI/WMwQTpGtu726DHcku7mHXYZaXNQMrt
aFqtVgGu172DKF2ZSkZ8cV6jcZGrTqfC5hMGyIPNCcfqUaqs3zH9qF+FN5Fa2fuqujT6czILeKt/
QEtaL8yHvEcxKTw/y3Zbq+I+/nnmI6iMoIaraO+DJ6Y+bZPX7UUoLQ4G+7UkrE+03Ih9+v9OMGfp
4wm+1f2Bn+j1AlKuqSQytP9pe6/3RbkWsAOj49+nGF4A77vIeHDvDJL/BJFnR5sT63zDXUF5mWmx
UJPzQ4/V8e3oDgasXeAqXVxlSVUWI8ymJjVelvixG1lshOm6flw0GS0dXi9I1aLB08aT0RQYdJq8
9n9xqHosiOvfeh8Pp8Et8d/rVL+ib2porOh+TX2mLHDvGvt2k4O3jB8GrDgL4zOTRCRcVyPHvfFb
YRMeD/q29vBI56cbzpApSF3HgfJfjigIUVYSP9v6wdNz+Fgw2O89/p3N+FwT2K93LOmpzHR4bVa6
i/+1qZXPKjH/cONvMET8+pKzkgFOKY0C7PVscCQqyIfTig1gBQtUNhDJVnAAUFqCHex0hrPrPveB
tneSmQ7PbnfTQsLTCyy+t4KzPQmktgH2lq+IVfCGyxjnkcjT/ZnLE4lKiYxkZVHTlo5vfnSQXKlG
GOjQQ7zA+nevrvVQVDtWh7EkNwYlXFWBMTkz2bT1XdozNoFy4Z8HnvW6B6vjCW3pRqFysqeZv66X
TtAgPUPCazyEB6QCKSUIRFbOY6ZVUuwJi2ZudSEcTs+p36bDwdjDvTA1MnPAz4uzDkNC/oFexBiS
+JBRQAIvYInElKNzwWwJZdzd5ZoUwd7dHoiUzKwJ6LGNWMxIh+8osf6KgeUryM7C2Glj2/72YL0e
bfBmQH5Y8B+kdEuqOhNzstLntsGdD6yDVIIV6p4UGD/ovCxtxSjBpwSrIXWuBIC6iJ1DsxJTBp/6
31/UuwpZkLr1Xjqe+Cxm49KBFZboh3uwEl1GNnKpGFTie0t3AUt88T538bMdbhTlguFZmfBOQsRe
EoasTwZSTJWdnwuAyt8Dvuvpuk1shQyKNcOzy0V6OA24eQ8vbN3vRblo4GLmmIvIt2z09/csl1aa
ytdUAtf8v5kXFWtFLmvIUK5tyL5YZAvmbBLqFSoUATtesyaKL53owacovI4hHlg7Qggi+XZ0Zej5
rOAqAWE/etbGoEc4hQ4Xre0+eoBlFPG6IE+v2Fegy4eVcoKKVUfD3czvj+qylS4yYgYS0eLIgcvm
OBRiCsoKeN57GB9HWYpcUzNU5CcJOrxdk5urJiNI22mL5YD8EUfFYJsMU4PDc1SVAm7pJ4596+c6
BL7xp/ORdHvoXQeVOkqOaQGwdBsmvTGuhUHR0FhJ13A5Ea4CZvO35eWCQdM7PoZnfTXDAsx4QKKL
uk9z97mNMHWPJeEx/Epay0/6MWAR5U50JjY6nI0zSrvsHSCsuC5vd0Rb5y6qFivfJUkI+ftU/Ywj
+5Vt321KJbgKAd4lTCtLSbUUNCgO81lWYjc5TRq/fO8aQSJInLPZpdJWAmXzWou64QQguQQhKJX9
y6TdpYggkJ0xxOAkMlxzBMD+2att1UO4Bamb0j8SgEs4Ng4xzFz9HOnsxPjGCkYTaBClAzj9xjGf
cyg0NrfWaMCjPtEl49rhxDZwseWY80lCPcVgwcZuvXZ4Wr9eSzRMF+BFynGPnl4rCeTU/gJ8TXD6
PAZdA+0yT/jDZ0KIufF2iwaRmeD/tK2y4LpsKAcX8EygSzQx/q/ZZb0Fz+MEmkeGljecDimMpxTz
54sjd/kDQg1VtqX/O0XsxJvnjx2BurScQgl/qOSsIFRyeNUalTt3xs1ApI1OseZ4I0JFVfb/gXnu
dBpgwAOZf1IvZv1ZeKM4j120VByw8On7g8xGtzrPt9dVw0ESb5znF8yNV8b1wObV+76bT0SSD9ue
rakzzJFFXZAUmLo7oEdNturAnv0hQnbyag3Q/jYrs31hy9cm4kaI1sFdA3YopduksNTW3ISnDhg/
UrQ+2o039/JcSp/WUX41johx71kDXkpCAVy9BNeRlLtdBC9AhpUCWOsijFHtxGFSWpruXFt0UuUq
8LrpnEn0ZhczjDnFOF9paKy93LI5fOiVYxKlRy8/gn1YRuWHQlvP3TAOHMCKpxU6BkhbfPBl2NqE
88fv0SjFFnHCz51gvztlAM2bp+VL/TTFpDAAeGRgIZ7+PfYdlZ28CFwaLp+kqh+sVUShTtqDvRGN
DwWh+ECXiaZGypMxHp3bw1vXJnA/KcDq7Br2TUNNB4LbOq8c4QkvMQ5L2s7uTkm/tTWpU0CEbHbj
PDy2o4hVULGsPS5qInQQSYDZS3wD+w87hC2iPLX+zk8J+7UH7gbrFGb+MPXxiHt8MNtM51qG/kzo
NiLXd9uBgm5F11ldBVxQjrax592U+X86O2hGxasd3dICbaqRaz1X4LqRbCDG83bzc+kuTvNtjVYL
gjFCUUt5M/Ys0bZ5EEeKsEiwJ3XlfupNbNu+4Mn0n3AMAvqiFJ/T0FoekZMe0BqULEzLfW6LomHu
3spZ0TiXKfrV2m8x+y+jHm+1fZCXmjStnFPTKQcXxa20JcA7XwnROMS1JDsdnpi2etO88O6+grZZ
3ndSAqs7nDt7ozJ3Vq9vQKmlKTis6A0DRvxn68lYJ8lZws2b3tUJIf1Gt+p2wS8Tlf7JflNO14Dc
Mn7gKA5G9rhUax643p8djLIV+ZDGQqf+ZNSGy4HceNqGoq84qZQItABMNozH4IL3783RD5CnRoTX
RNmOD56suF+Jq9b4HBm3Vu/79ASBpL2eg0b+nNuY/5Kiw4/q2pxRAPMhDUS0Drj8GYtxFoRj+S2W
HILuRNM9QvwaAnpa4H7V3sO64aMpMi0CpsArk1imo9YNFCs1MtSEANrwihDhsU95hssNOG3E3UT8
rz2XXsxU5WSoO3AQLgqL9DD+nOGE924aiaQJS1ItVpuaEHtyyoGLLzVqTeLv4CTXeoxKct9zNtKT
FyfW1wcv+AokiOyBGwqANHd8i47lNL1x2CcTEPj+HWQldZFlNCxpx7LGvZS1iAm2KlOL/haVfwoa
jZd935JstURQuTOAOJ4cuaHmZfJQ79QqWAjt6DU35ARDjjbSkk+dPprFZwd8+YqdBPzkTVJJetUz
PoXbW2IyuCHARYasT3VqCJh/wIIDlRSxpnZtCuX+Fm3M+WbEGXvrV66A3Rdni916/NKuBs9j76n5
O7IL0CCg8wgq8BERZoIcqd+aRIWQQJtmsn6iqjcCdy/wZKgA9Lbn4ASuspIk7+9V8SnE94aH/fF0
ZNHPl2bbYQHSDKFw9rHOP01b2CVR0XuhS7rlJgHNsNFaF3gE2kW/irlvq+b79VYUlz9yx3UTAl7z
npFqfzuE0D7OnySpVAr1awAF3f390G4okGJUKr1taq0rRZKwr3143SVdKuiDJ17tO5QaicmOVmm7
JaW7UWmxabHl7sy4m1CXFPvDR6QJBu7MIiinJZl/mXUYfumlmC8P4XOB12kuWPdGYIOS6MPg1sT3
3W3Jr8z0lNcpHYpDSgHWJo0hRXjRgLbS7LJRx96VcPtyGeOl+AwEH74iovTjuy/wLQ+NeobNIqsy
7Ty199t+sgXT5dmVaMUHt2BaiYrhjr6o+SiY4QPSj1NRJAS0selxA0sygR7uUusz6VHUvpl/cb5d
3UBt3Jns4zTCb71Q16CX9WTNiYn1uWyup5B7bExSsI+thpf2hCJ8CO3NzA+wwmPHaM3c1kg9llyo
tFTdCZrD/e5575mIFJkRRghTvExCa8LQaTpqdUENp40g40EH3CGSQUPR0pQRc3IS790Qc6dutB9a
fjdmjh1rQiGvpCz6EV5MxksFvrmQq8IElpI7X4Scqx7O1ymaLA239SLiRnPTzSnE8GIXLDDPq3zl
joK7bBMzM+26V9h46kZzMMwisjqO2og0byR+rtac++hwsRslbJ4DdaSEwY6bQXEfksMiiNUtZC+u
46++/82CRhgS7mFMN+yv6o0JC2lPbcxdEbY+Zhf1b2LXreubH99l6Lzo+0VKCl+DZpKMw53Nzybh
z0ZpxC2MGAupz0Fv22leOcj48BUpHfcuLsxpPd0x/9sB2teTbY6tKxoLUDvd74/erM631TQwTMfc
qixrkhBqQa8R1uwHtiNt1oz0R/Mpjcd84M+POlDBh4uKPY3XXxSVwA/gQKK8EAbhPhIQM0d0uU96
P/zpoi2kz5JTblNerjTXBG9vB1n0ZeCgxtDN3Op/SgKllcjbhBLQlnlkbICgImN79QPfl6KSVT+E
l6wZ8JD3pmdDqI3tUB35jlEaKijrzD44GIcBwL/dh+SqxvuVDAw+69MLyc80yH+A1ZMBc3hANENi
mGhN0K/RjK1SsrAVuwXPxz7/HI2eW93m/1CiX7tjF9OYUYKbNHdBRVilJsNPWqSSCbHCjSLmtkrE
RsEkj57bmSg8WzA8XlgSgQ6VyonjhH/nWQQ+/x0bpQT+1ni+aj8MAIxnVmFBGeIBsw/q7040I7VT
SQy3YeVql0ylWnYV+JV8RPJPr2sVoH5btnuusASq8wjF7V6P4S/z+JnjmEasskFE3OwJeQb/eXU3
yXPnGf0/oC38GCETGyXYJJmQmfBgUlynfuuYhqUOuQrtL7xSbzc17BwvLD4ZB13sCaBm1xQSBn3n
67bAgV9iWbAgytGlrako94/B6mVze588iL+HhsoSQZhHJ4eX9REr6ecWOsg6rg0j00gZezurlotE
selfK/Mro1Wo9ubrmv0B8YrViyEtFiSMXc5lEfYL8opV/UZs5A7Cr/8gfpj3FXpqJBjumyICx+Gl
wRqSJdGukXaGVSrx5oq67vG473jbtrC70kobr+OgTFprY11krTxwXuy/0rFodF35a1XDmTGw2gx9
LDX5fFos15dB8GfSgzBTeiaopdZS9zOfEY0AfodkibXG1NSZTmwGzcAhkAc/TwYUwjmonVvbr9X3
PDz5jTBGtrI19fzQuN9e8GJ8dqanQkQuJJpmQT3+SMMe/pFcsbTidm3bm1RhykmWE+SclAYDXPwW
TwfI01ZGDB87TL+x9diJgs/UxdpeKSp8RLrEzSXATMvFV6m4Bb5nBXLzTIMt8iCRJvUPphNkIwyr
gvClcl2dyh/tKf9SjO+K3omU621HPOQGFWGzD/TgytkZNXBYjTDlsACaoM+2SxerkLKLK/JXndtY
+t4T/8tmzxbcWiW3jma18EkkxhMsmN9ce7dNpIu7WbqrQ8FjUTW+bIb3CFDbECBFq14V+0QrulVQ
KVFhifs36NnhLnwWW7v3g0WuauSP/+Z9jLEkR0UIgCmuvegouknLtNeS8BEyFrj8MFRHr5vHDFV7
ESYz6XTPYzzLxAW/rSqGPFAhqnajzONUK3BWoeZamcs8DuavrxbIe37Gtx7mC83TsYUG60ZdpWcj
aANpWu9y81XIKBaKWjsHhTxy8ddHltC5YDHuo3VgOd2afpxO6209iRHkNBr6KjgRxP1Qo4kdzzx2
KWa4V7sUQJa840a2X0GTZCqXSvbT5rg02a5BvIgD/f5G4DwlpoQ6TfO9VOht6bPAH0NXlpeyDSk9
k809R9oo+7cFRD6vVjStxMuWWtX+DMBkPaNoY9ZsWqrMpNcvs8BBLAnf2rgCRmhv6XJ8yPT7/LnU
HTN5iqxdmWYDeJLJcJOSoC3coEyX8Zx+R9az2fITwp+3vl5Qqhdymv+As7HudHAWesrHhlqE+827
W9mepNFpRbjn/MBchHqh1FQoy/Y0XhLP+3cwhCTVa+HUO1YsvnrS2PilUaOMYNDe83mcyGL6Rm0Y
a1ZGQDK4PR2nPKld3yrqE7aoxJfhJNkLQSkHJghJYazUC6Z7i3VfE3dWa9u+v6mk2t4vndmuvcYf
0onrtfQohAWPYTMJ2yVozZeS+WoUTybTfQpNNoLY2gqGv5VO9TPhNy9lepCaySnfh/T8otOoSC5n
T9UTdy4B+1B9FiRxgrIufZdJL/pV5AueZfjRtGB7guk2xThY/FhNba4rjRTe1wivCwrhqZfqrdhW
u1vBPcEWDhxFH7cuWUn49kGEoC2h4r5vRwfcgA+EM4tLHpTxg3Z94rvOovRjvHDSIshslyZlpyCN
02JHQzh17zJHJmsVvSISMto6H/m05U+lf1amg3ft3VUWl6/lhc0zVgUW2FxW/9ORGDTRELxsnqjc
flOC3dCviHa0/23tMazSFP7fv5EccZmhTissKUkJ5sqvnrm38RHYwlxSTkhlvhqhLEqSecWpTnl6
TDzNp9l9Oj6yNxw40PrrnaLMEcmiaQxpKLFr8kXoAs74sXu/mFM4YeKbp1Z4hg/8dV9TNjM7AW/t
f91o0mJ3v8W3FPCiG1s72DgeBOJPmnpK6/sl5JSRyYvaROrZR2EjzSZnKdAQVWEQkD2UEHt/DP6I
sO2E10vzAjUu0YxTnSd72MkFlVKsUVbA9IBad8dDIv1fIIakG+r0/OEUxYgIU3CVm/ZqBMboY/6K
d7tTcRYkrmEDJAYgVj2ma9qeM4jL7syk8AX+1gAdCKErsYJ05cxDFVPBERDDkNzXbKklh8i/q50s
0Fl8Vn3PsZ8C3dB415eoz0qrQ/irQiaYwsOjytqTvhotkDApwO/MLb3Ly9s+bTd8ulum7bR4lUxF
mxO2alTuWGMqhGUbGV2bpVz9KHpjb2ZSe0RE/ycMj8Nc0xPNnqxKnVCGN7/zzLZHWt5FCDCoGLOT
3DJoq7k88fTniihE+IVHHF1OPoYaPVa32VCc73v0Kq3PWVcdn/VE4WesPd89/h84ZsgKvy3e6jQI
nKYqOBMhTFyyRWgycPPZPSNEs2nTGjaCsZLyub8ybFYWtKy61Gtip9+4CIevLdyx5Uxfdjslt+mz
fjkKSY46qc1tbBlnq3TqgCSnFNGnw2RZrUt5SfX4qD4c5AOCdhIQ0rmIn5k5Wp5KqYMolYq61Gdj
KsZj0VzHVqWwhKsKukacIVpu9o4Is6LU4v8bctdowoIG5XG8KtyYhfDAf0oUoLF0k93pFg3FcHOu
TBpSs8Ey+JAdKavVqprxqJMpMl1jqsiS2QcYPzniKHEuVdEm3tNrpg1bqn4IRaTZBwnp0ZI9i5mO
viz1BwrV6j0L5ibamLzt12lnyU4MtNUQlw20JFlSKVZ5t2FPtYBIW9xNiULROw4E8Smrpy8mJfDN
l6nAn+6kC9mWQb1zSMVA4kk+GpfPVqHeESCZ7faTjmZh33uSWkl3foOuczR18NPZ0LhKnH/94it/
V69iTgJAo/GQu3fqystuBXUMWUz+OdgD/AJ/WYms2blCBo0mCjNYtXYH+eNIru30XTiI+usa48ps
A2lLGYr4scsyOlcgmAKfeqWoTnjlN1O7ZAa8w/iDbXwJserw2nuhpKuLzppK+cZvKlenQ9ngdvb3
M+cIWYNOkyPmaLlHdqyDglbnxeiKy6EwtUivKSkDaRQuoTHDs7r9azLZl/29/Tj9BkkAZ8qTuo/2
CkervhyRxPE2BsizePlK965dzJbk1Z8pTP+aHUAPWe8CCv9nsEBQyzweMWFP8ra2YLpHPTANrvrE
5srkqEi4bGX23JTUvG8eGtaSwXnEeVaC1A1l5Hj5ZVk6hudMuMbuPFDYjjfJgOW1bsbn2PUr41b4
TrotvTCLw9aA6oyEMR3zab0diMUraY7W041pLRzc/TzgkqMiujjLFvWYqE8Do9GsxyFAbYqWvipO
MEsjsOAg8Cojcj3lLaROqpVlQEQLCzqpfdvvLkfuKmds7L6IIKrv3T5jAhuySlTlIG20fzDKb8SD
redMm8QG4fzADreKNon+Nunj5nOWdZlQFbx/+EAWgX+MQ1lpKcwB8kujsr54QDDdOrAV4GR3TZbY
1oFpbZplmLmK/oYxRIGJXSBUOohD8ji1CMEqWJ3BysneIExy6vwiQ0rmDsvZQxIaKYqXwAuyK4+G
x/Cc765awPNWJmFLA8+CPj0rISKPm+kG9kSzUhWSOG3OjBEZ+iZvw9Urp8rbQnUhi2Fjgj25rSuq
Pz1v9jSSffNy4negjIrGewTTADSEk5O62kh1pSCUvmmSUsuwUSNvwEVZGM7VlY884D/3zkKrGGvo
pgBqT2LLVBET2BxXe7AP5+8ni5x6+pcjcrjV77/ci1apDglfgn2yDEqMTXZ/iL1WvnPxiElUzKkW
IUVX9hEY9D3d847MjmuuHqhGz4DszkGZs7vMzr25pf1zfuETGvtYlLQbt0atkRiEfp6zrz1YrQaq
EnQdLlDhDu4mxizFrAu8rDgs4MJo2NNL00CzR/gOlnaEUeVoVR21o7lEISA7C6tdgM4pyje9tEzG
X/8JSLsTTKcrMlo4k8AFyKFJkvi37OX9Lbut4+dSQ8SNg1DP1LDT/HhT2P7313OdJ6vfO1mKNtw8
noMF7QP2qt1UuD3XLtTjGDsPzXwmSB0YzBjXefPJe/OrK5zE6kRgNOlIYykqcHgPPR3Djs7r0acU
BiN5BH617jI+QLIPgfjAQjH8R/pUUc3FZoWQyTgAOM7BkowuSls2F+rCKT6AzfMPufYI/AU8h2go
W6uD0+Bt3tk/OGXaW1+psWB1fb/AE+jdnVi/lG7sJCscCmKHldBIuYCWFBW164HWMLG6pexPdIBo
y0rERs/asEHFlo35e+2xwQC1rPRV8vAGulImgzTud/TT7EKfkOcvmd8aBUWyKPu20/NGBSRMcCy8
b29dmRw75zn5RElinXak/R6ynhrKEowHDX9/pZ17Dfy/fAMw9ccinr4AoT/DTb81kD/z1fXYhlcO
G/F47JRmGk7Lzme0zz9qEWcci/U/de+jPgIba7hSblhupEf6CZ0SZ/e8oKozMn1R1bt7nl9xbDwd
03Tgl8jha2CTMbqmCgTcRIvJUmMegCBIcKT5czeoNV+eaO6hhCSq9ppEvb5G5UEnx1zSpIL6TnzM
jeNDYe3xQR4ZVxycur40duHg+ppK3+i8HP0RxFeWzYwvHglWDq+kEjHCoEo7W91/NMHG5XShmNK5
UbIH7+1TTZW/LU6oElWGqXkHfx6uNGhmpZpYs5blpkQAOyDOPyo1NP5hVwh8nsEc+qzNFjQhPIZb
+PGvHmrpwYKVIUIK9+FHukfBA3RI7Wx6Dy01lKSr4cgntWyb/iva/IwBo/zvupYwfUtg0QF9DAkM
Izfq3Lx1I83SYNf9NT4/DirvRqcakUtNucmFp6IruD3gyU7Q82JQlvw8N1Al2YMVzPAZwkC8pOfv
P4eVANPhXQvuFOk8iht/qE2JZwX5xPoTnpReM2UNE0YWUU2GIjgVUuutYX2buZronkjfDDOBMESr
Tt9wVjmpMpVhDFIp5pre9faj589AKodYo95v4oMH5w6cTR86mD2xuZasbCdiqrvlMg/Bl7h//T4+
KJd/g566Qk1NKxMlgaOK1E42dbTEWHp/jos3FBGHc2SwN0oVj4wQ8ZgMX/mJwy4yHNpGtFsULk+Q
ynHVjEmR/jQf/hZ2x2R4wNm7hRu3wzu6rqKd4bwr6T+zi3J1tpR2Zb78nDDUCwSL013icfDqCETo
xqLqw1djcs13rIjs8voCWl2qQLW2fmP6z0l0o6DLFGAW33w9hWs4jtD7aRrBS4iM/jAmBYPt3cXm
GiZsIaaSQLHPnOdcovqm3FebplTSPPy5cl7laewZJgLHXqnLJYVjHGavs2Wpd4R87nsTwoY74U3m
JvBVO0pmsJ6RE1rdcK0ZqYkU9O6NF1pNmPWHsy+XgNn05j3wzrn3GhQfI5x66TrMyFfoH7rMreG9
5916fLr2lR6Q2L/Ts9HK0B5/GmZVh7anCX2vQ6RFEWjvqstmQKp/2o4l+iwPLbIH0mNkek2PXlvx
HxLFk4IEGvK9RxBjsd/UNazHztPNw7Q0ACZP15jk0DWwZkRxUEwjzT7gVFwlaICT3LsHREh3cA3l
pBV522koNZh/C9smD8Sl/jbsmnANUteuF0K3/rgnjAAOF7+nhkezM3rxyoEH45NzNQqwkoSC7gsk
F0qdp4l86IvrSalFQ0Tf1DG9kKRpbk4C6WA6fEIRUEsI6LlfTu/xxOLi/iIP7W/ZQLq19p5aNq6Q
d12h0G3mOvDyMB3oI3a3PQSpE6ot727ur5lOnWuR70jriWelVB7P5jta0EVPibbxP26XemyJm0yr
h31vXSvX3SUfhsk/Equ2eOn+SJG6KQH4bJL3a50d1m6yJCqTu0r1zuFPq+jrppQr1snd9VK9BrOg
tmipZ/sSmYTulGGxUT79kkOJqjX1GxxsH+ue0mga1ito3zjJN3bt7lxZA9A8YfYjEgVM9bSvvj6M
EWO/nuEoVpv1ExvZzLp7883QpdzCz8a2LuUYd/cZ2DFSD9sEW2uUm44x1F/6phXHvvsG+bluVjXt
BoCdY1NAfRQreyz32Nq9xa8K/J9jxdjuy3pSXNa+fQ+PlwWNSiGdXqaJv8OZqlM5zX3EYJ3r2ymM
FUXQjqQoImWhFojAHOxQ5we3ZOoAttLjv82muC5V0oNavUWiWUgQTy95wO9NbbtpRQTmzc5sdoM3
vmtIg+AXl6MR2Qo10ukJe+2Gv89xtLHdVWANF9CusKQaqNnWAZeMD7tWClF6JYev7ORMCaMFtIsa
RD2oq0DyVvNY70wA1MXGYLpWgXlPv11HoC+78xFZj3Fk5saDcjla6Xv4Fm9tGZnhMqQ8/GGYK/8K
JYvglothJyGQ+sEc2y+PskL1keuupL9zLyAR0FAKYd2P0ho/HU5AEvc3tMtflO0/DUwJ4uvX4E5r
/EZauoqNlhwotCfg1BEA9hgUSWRX2Mxagd9oXo7a9uiu8R3h1gbK1aVvEUsM4uATdVCugznBWgAx
O7qoebesvSdqPtWxqKHIFxHoqQ81mwff6h5Sx47LJW6+Ga+VATvIhCl0HkJtKY9XTd+zn6G3qvSP
py4LUvY8ncZO+jq38G+Bpo3pf8lrI3rj5mXixQ32hS7sScnEGYZBjJ/uspMPJ0LQdrID2MQ8izH7
HJSxJhnQik53P6wNzn0Gpb4tY3cuGb/oLzEnImU0TVqGc/7XP+yru59cksSshaQp8sDxBC42jZwx
cQQ2iSaydbL3BaBwgd1SyAtBGeSrRUrkRylKcYTa/2j2jag4ZylWDZf4MyRzGcuUGge3dNnFZPYV
gaandHK6As7xvXaWVBVlwIpXmWqkM8zK5WmUFnuAKaOwDMYssGiqLyFQ5kztgegzHOxfImyf2oM2
zTagXmHr/5JhDaS9e6/KTtAqkOv6HOBM9KhE0uMg827MvBezAaVM48Jfij62XDc1+kPTaPYepy1W
lpWHmVL3982Lgen8K1HxokvrlDquNfdY8XR5VljHPnhDv69D86dCB7kPqr9C55byY5wp8NZGS8C3
w6F+Dne4g7Ci+XbYS73DmmSGuG209hzHznerlgfNe1vKXUM8dBtmj+T6a7jO1XqEyY8OHoKi9lSA
462Z2+zpRWFj9AufBPfohbLnNSCT6bU5BftoKimIWxJX4MGeVwLpjzvb4xqJDAl8pAd1/uL+/UnQ
FCG6f4eQnR+4JBbtENx2hr5LtzYdoLntu2XYcE+IJUAkTIgiWL3eGEcfeHexb4aI3iwKwayl46Lg
H4Uv3vLe8v7SZLs7Dq/70pYPknvIo6VuDG6k8xAkWif87Bb1rAwa0J7vWJuaqZCCPhMPYNXWsz5H
OAb5/HQ0IsrbK4kyGJrj9a6Ee5HzkbQn5k5wu8xvI10ycJHvKkrRkVonEEnm6/nhgojEcbKhyJqR
HUGpTnbh5Zez5DH7nyohtBePcBN3X4vYRq8bQSnrJ5leuGnaFDV04V5T9J9MQRdSFfqBg+sJG49o
yaffKJ5NmRglV0uZldiYrxSZheQWNuatjdaKR35lT3TxpC9noRa5XI3Ym5f4hZOK9ZFt8VLzWTOy
9o5e57SMs+hspCs9JZX0cjk+seT/X9PEaAbLg94oa5Z6l78euNoTU0dfJE3BslMC47iYvhsj4hj1
7umOehpdllYn/cOvj/MiZNWRyfkBlYHOQWtaDnD903kUsvIjANPhltZOHQrsBoG0bDNNGOmZrvR4
An5Zs9AXLsxgKmz+BM19ScAuZRZPPdEllaVqtVodMbJWKLYsA8OQMqjQaLr8QRpCAxbyPZT4tkq5
LQyw+O8ry3QT2/m55lMwoIo5XyLzh0u6/1mNbBYqtVvDM0Dv7II6TyCdXZ79H3eFhkfy2AT9PjRz
Joiee6gmMMgvS1ljnpyeJ9aLAD17hFKzDpTew14ZHJJQGACcwMPp29Lk/TtD4EjNKUSvFWQvkKzt
qIDSxXSKWM41HegP7EWDSU5e741bjQJTUWa7RT/K34mQ49uHm2IQbT4mFdbZEyD02mSReGdmH3sv
5Zm1/NP10MsRWnP2l2YTAQsxYFnBnORprp/y53+9vRHtRDn9Cesc2KPk524eUd0FuGbSKkOr+w0G
y3g/iKtn49PNwM2FIkbzBvJ2A3xyJk6lGiaXe9s5RE01aEXhSEm/QvMHE7XKECFzwoFAmGGHUx2T
+I/WCPgrf+SbBsgu8xPPAUkVIzQ46apg0LzOkTAxvvTxNW7A8ksGHg6YCudZ3s++u+anB9yGVnF8
IKO+iLSznGG91rqReLo9Z0XtUPFKphgih5TnTrmzvbugVwiynKD+GqtUr1Avpz8mQmNOcSGk21ht
YTYhWtuIqO5MBIrO0eCT4MWlkqLxohpUIxfACNgSdBz10ihfM+WT8anJ43LdmhyCtgeeQ1FzbRuA
yXdFlT7YOTTM5CMxbkLcy8d68V5FF5ESJwCp+zn1cpLQExwSoPgZurvOlXvRF5+9U7hm/T03/5Ru
zW55aP/XXXlF5MEgGIgXPqILM4hvBkPPpaM7FgGD2bCK7Mm0sD3I9nhaMcxBBBoKzg6iJWlMtvKN
fgyFokMPPhmzkrl0BOuey7DVTFLcxeeANGNdLRgjsoAObOad2cSBu5wML9oGBrlPXbjdF6K8HQaS
BgHkm/3o2PPlqcWnRtq0ETSMvL3zwbW3SNQ5KPZf/phzW4Ynpl9toVZT6C0kQwrKnpjDWhC46Lu/
kKnuv0na13b/pAiAFHJySlcN2RBgLHNsa3jQoqQ5qzuwzuA5A4Yw5dW9ChTjZzZltOFxXxQWTAJY
OKisd5YWaQKZaUkjEQIYy+0a5RUiO863IsXIGO2QD0xIMpJb5Wcld/4Qn4NW/77r4x1qr/GRVCJC
qR1Pxojk2cksNu8/gHCctb1+0Wnl2RwwZz1B7cvw9ggv+w5RN+b/oAiKIsqVaD1bFEL7CYMVoELa
aduqnoRrztscbEP/vi8Ty84Q55B9mUCIqf+JtX4vmdkUnKfzJa9FX9+h9HHzhhkbBu9NCWUkuIrW
pqDM9D+oh/508SMsRKYPAYvUt5bMcB8l+fBi4QeWs3M7MWobwPWcM/1Br+MLWo1P8rlF7xt/BOU5
xVibaJI7t6WGYGpylqoby7B9AZ3iq84GWaOh2F7DFf7CUGWKJclQxTdwmU9gCusnXf71apHFcnQU
r5IA/2LmWRUjutFO9CbYPINOZALG0tLBDIJR/sN13cZGbzZ7Oeh9zwDw6WvMKnFo3ZPhIpjqGliI
szmGRcpS/j6YZ+fezH9XA+143ppLMkV1dD3X1izy8YG1neFv6RWhv91JD6FTlKmfLT0LzIQukm4O
C9ytyjNVsxG5tEkE1zoID0n80/pKknz8QfB+/VXmOvtt4vZiNt/de316p4xw/SOMU8xD25wCv6QM
0CgX6Vs0zmRFcVlTPpNz1lPXq7MtjUNvJ5xh+idYOf+2Qs0wWSyUbsR2ERjoo08Oaghpijxr2SYE
xUazkqY+8ImpGzYtsIlgcL/P5Dh2hkpDjgokykkT0U8e2vwDpNm5PU6FpIVdmiqfh0sHu82s5BlG
NAxmtZrsfy+tguoj/UsE8F1pvkoXvbpn8DOEUlH2oiDpKxQ+4wAgpELxPfiWwysIiDuvmoc6101T
Dh8FbH6o5IjetNhh1k0DvmCJVdWpEMbWar8h5A9z/Spuuqt9yDm5Z4ATW8ryDBgvx9GkVfYZNhCT
56DJTfLD2/mNG7zdEMmR5Ys6qUs2dP56gzzCgWza2jDnRKC/8BcSsfHqWrAbCmxJFnoM0LQtfnlo
qJ3iUsC2RTQMzAGGvbliRDodyrbPy79jFOsvhXWbpiFenT+4MX/lytN+IKoAS2qLjeKYE+KB2+zu
ZyafwikXsi7SgmYUcDWF0AteaTWrLk1vNX7hHtgyXYOtsFtAAOv0NCN8qAahJipI2hCsvEQ3dU57
RudVugGhQB4ir8hhYsfRM8Qh30QWCLYIrNzxd5GnnsiS4erHR0zyr4TQ6Nnu30xvVlYBD+BslUBN
9aWKQPPe7gp3FLxNElZjJA9tjXLASktqUF30dlJN4C5dsDXez/ED3v+2qjOTq26fQPdNlJdBZtx3
rjNexRiGP2p7aztyCGzQ9VIb6LJV6+OvXKspffGB0b9SV/4zijnPYDAHZ1lw31IwBrTeIqjWRuV2
TmfrWfiruLV06/liOiQDSBdU2AifeuMl7gmXLjPp80vyXKMI1fiDUf7BONHA+a4z5/mHp4moVHp5
5fDQYfQyKiB/Qf6NhObPg+4PdWNABLkHKKVTLbvk375D59dXTFtzVMxfCACPIYKz/8d0iIG4Q+f3
ABBqOjeuU+zMP0wrt4KHU8AgzNjYE5RByNKNvNXeMIetTTRQSZQr5rXIzRhN1Um8fqDl8VyIROvH
DZF3X79jSiSzPoASx/Vbg01aaNQ4z+pbtQIgjs/IxPskdk8HnE56rXPEbny6RKhXW9iaF22IHutb
qRt2b/V6z6DSh51SIrFw4KSCIt5yIxlxJGjjiCIh39utUSs+0lLrNRg/XWLoIIKjqw/7xhf9xOov
3IAr8/QCW/wgJVNZzhylWqD8N2xHWSOkyCqRlVeCHSYN8+sscpGAaLJuTE/LO3EVQjGWHw8eQAWH
PqJ9OXwzM8FYD0P+M/mgFAgCiIRAlEEPjYx15Te8eZsi/ojoE+fNTqK02AEqlLIIek1etTQoo/Ww
mlwKvN6JzAwisQPWaIFV50Fs8nERMj0RSg8xcrqsmd2KqF0vHTlDLOLox4tR2mj0ITxoNSH+IqWs
OUptn5FSlpxYFh8dLxEB2ua4viyu5b3cwJXr5Zqgx+7K6/Sq2k/0d/m9KROCO+wAzDZsB5qa6I4X
c3hpEO84ur2C7CA9dbPI8r9vkfk2Ts8QZjKZ1e8ASpcOhtC7YYy/Ju5Uupv5hb+M2nz3GwujlzQA
0wQa8yK+ef1YyXhjH3smBWs2K3UfpjUOLbf1l49c3ojCMOOj4g/754pEBswf07dqLM1OQui7opSE
Wp6wUCdXuxNZUu8eFGmRWAH/UeipnEjexPuSiNgHKi9L9cqgt0vmOS0X6ZNzeSevTy7BKdrR+bVP
9nkOGd5kWeE+Fa+oKBdZsm28gEqQ6N7oXQPYz1gFzLQex0/kaoAO4A5z+kwdX/G3+dfSE2A6IQTd
GVERv/QlNlGXcsBFhQSIZSdwQmMWHHPjJdEU/koypYJLVdayrP4UcpkyszrZczuba3yih0VjqxdY
aTm58+LyR75hKmc8/33sVy/KXfbEEqfbu6cFyPxIwr2HJgsRzAJe7Ym9BBv6EnpgTOfQtYAGa0qh
RcvWitNiCMjOslLUT4hvvW20skGMUC+z010MAbGLz1L1IpGac2h72jc5XGQwiGnkzvREtpwY+IYe
qHqCfjK0HJGSaVMtrVdvpHJ9EIqbFaeLQapEYyXQq3P2XfXu7rXzRbI21Mptz8ahIeQIgHMXfUm7
1JH90yvbx6BUNXhzXqpcDoEfF2P04VL64J482MPZo07aYKDHFnceROeCjYnZgw5kJPOf1ZYXr6IJ
+BqCiKlBFGmvPmfdbpGJfDlzBRLkEj+s0ucHE+S6K6l9Ntd7J/4tR5VZQFuIqIdZk+obV2zqQs4j
kI/eazc0M3JXemEePbE9YCmY2P9P1+9iNrbdlmYJVJ7v6SmnV5LnEc3IEKWR0eH78WeqKfob4lIw
HgvNs2DImrzETcUmtdTz0uzhq2hbXaNkInAcUk8LFHn0p57pFfw4C7Usdd+/d038M9BA0/D4RhNJ
Vd3CcPmsk2+PpmGoHwTBz49J046jRQxI4QiiEjAUWsdNLCPLvRt4QgIpF5JUNKAe1+mByXjksd7A
FNNPOF3NHDhPm6K+bVYTw/Ge7LwwNrZfNGoLYZFi0d0ACPDI1rlAQPE4TNgQvkcSstvN1IIib/3M
LE6k6oFLK0ci4P3SAChKjlFFYwlIzdYt2bxkXCYPsnE9x5RifF6Z5KB3eMJB0EUa6Le/AEJTwZHH
2cEdjntrxp7weAUPrl+ubCONb5v0h7Wki6j8E8rmOM2+NgXP6GT4WMBU/26kLmzhWz/YymbNl6xo
1CwP7dy+wAKQ0ThndR5IsfnJHFD0bIlJg/DueHNEaJME89fhwgfUoU2yzgPa78yVnNQhOAsF9NOT
53d0RLoAIxDoVkxVqELtDZdMF9M2csVo2QM3YJw+wa54Muyt8lYmSlZAn/bzOPPlmryBIzG1DTsx
uovU2sXWY+UcXlD6XKqIMfYYFrF/wmgKlRaWsvPybvwVsjj9VEiUBJsdT8gfhhjIqK1mbYbmBv1s
20SIN0cAx0eDMHMTjHWk80hHsCsc/wFWH6rPaeZpRuP4xFRY7NNBNArC7mGJUP+IXeBjR8bx7uyh
u6ioIIsyrJ4nSekyd3GCPCOWub9flx67ZkB3UHIL3lVypVsqTsfV6yn5gW1aOwDjWZ/8zKM6KR0N
e+D1uzhgNBkox4pefIsu1+6+CkwyMfl6D8I6xtNOAN7C4AU8k54kg1q7knOEm7hNZ8j78Fob0pDW
/Ay3WQzsxMl04/cqwQnjCGGiukdMcrWCQCEka9DhDmAb5c6yiHj5c9XTzFdzX6p2vDR3lrJSgqdb
LKfBmYlnvuTu6zifzSPO88seEjIKwwCMNpT9dwZS0aZQHZVLY/yT+6kcA58wMO54wLmsQ6Tsgrxt
QPWxquqCwM9EZ6ChlzS2Z5zLXF+qNunrd2rnXno8XF7JopLX9qSRH6NfQP5W8MYYCJlZW1RxVg1q
ioZYi3kWkWE72GjUQoTomXd0r/uWt7G+Q3htKUQTg2DLeGwiN9CW0CCIEcO6ZmMGfC6oJRsFKvXp
OiFwtOOsWAb/JJLATkUMx3eHbF3vmxxR7JgM1SeoqJkccw2AGZrPa9T1J/PV/547RGLB3kIvR5qb
HbUICOulMLl+V5Cbzb35Q1/WCKW7qyVmXeHXTcVcq0dE2pNnnycdfOLsfAyeaSMeBBJwZsAJP0oU
NgUF0bCcNpdYr0AoxkJ/nX07F23rif8cAFHCpjzLcpKcptZDpvqezheCB2DQFjPjake5kU0mSe0H
bhYpF6Hnodt6Q/GS+6xdfss1SpREyG6TYnyPLK+C3gNY0B7mCqr4R6QGqKbE+ZHRpxX3BUln5qCu
enCfdKYGEWYq+Bf4PqNzSDJ4B7l1YRHbjJlNvDe0voiJ2l8GJmjKh87STSQKW65XWEu+z0oDmLBp
9MB/lFlNXg5yh+x9NhDiqec1E9hqOmmMltcBbzb3nx5JsdzkPRKCzu3QDqrTClkomwDBCAFU0QbO
cd04FaXh2m5ivUfBBbTv58RwWCzCvruZ8O/eeF/4xiQNNoq+uqdyISncjglyMOGFi3uK2FWfhB/I
1vCy351lLaguoxtqnRyBp1pOnjZrgSSJ73lBez9ji8moe3dr0n4LUtnFDi0QaYmZYDTVYVAMhSOF
i+FB4p+57QGybTz3NZNfsP2aK0gFL7my42bi6hWMKNCOZIw8TCekuSts5Fg88pTdrHCc7SZUxGEM
PJSBkPhN/faNIfLEDV4b5Jl6irxg1BcXL5CEKdNcV9E9t+KFSlhizGNpO74yDVprynddLFX0CFCS
kJciNl2gibfcrmkPRtlpvWsFdyqnqrs8+wl+V2aYpWw0/toPNQfz14Hw7Y7ystTmpAqhnhaxYoYS
6l9IFwObXgSgd7SUvsoauXbmmkarUOGNCy3B9c2VCdwDja3L+UuhTp9m0kvT6Z+Hukye9f7FIW7o
097ghHfCY20tCMnGGgyZUQe3j571nfxagjGQj55NXiu8Ss+YN+mg3mVl06nc7oKm0jE3/OVA8LYW
ZGywD7IxGG4vByvb4aa8Od3hIsxkbgj9wxyl7BqTH619LH6YjSeZcxNroqWGK9Zj8ODsXcYIfMSQ
fMho53yvGTR50dvDRRTmkgqGybX77eswyUjrn+sIATrAgoRyuQSXRLUoGq2dBsqcl6EjDvbiCZmK
0kQaFdrWhXH3WidrbSm+4LNcfVC3y2OrQ5XR9UCAZfCjqUdQEvb7/52rbqb0BwbI7TaoJqzB3Mo6
/KrWp4T8A9B2PtIdHEM0Q4yY+QfwqICNGYt9ovZR0IdM920Nv1Wf6Eyhd2AuG+BvYkHAJfiYAAyz
48qjlZDyBoWk03nYj5zFEBw7E7HoXqBDoEbN6XqCrHq8Dh9c/Fz9g9nZhIvCYxNoB713d97am2Wu
PlsOnj6yWNLZ0R7aPbDJkxV0pDAuDxq+Exlj5FTupKkiTWm2eP5LTf3S2Ie0L7oNk5wjWHmiy7pt
nQsqrzHOBVQyNnE7MlVRS9hAAPS2uafvZLq+rPs1YeqZxN2+j+ReKp9dNsSpDY6LBVYN1jMRxVRA
7s4MEVXVuOW/8ZziEz2SOF4p+TpLdObFvBqEDrIEA3E2+ofRufIw6mpXg/o2XGAnEUZGr+4Cb2nq
rk2ykJqhhb0QGuucSjDfUM6Kh9Y4aB8rmfJIZs77xKPbd3jTlyVROxc75KGW4N1QOiYXu19WM5U8
NsxxCEUIZYkCtRN7SCZ6Um9AkYp8pHIlP7xhYnd/IFNUI8QlDS+Qt4dAjhVCdAW0bk5GRda59/J5
Z8RwSWnoPhqUnbZWRtbe1UlQRAaZ8pIJgisHR4U06ohwC866WD1Dhbx70i84B4+Wvdt6SPF/j9fE
VW3huEg6kb0/KF1arrH5icyCByl6qZoh0egfbWcB2PNTdz3n3jieTaZDkaEM6dMQA8m0WL3TX14O
X/D5Bo/ngi2FPjpntzB3RNc2YbhX+2/anQbfqUOHdL1wt06H+FC39D/upYLXvq4cnyqf0lE3A338
C5IAF4Z8hy2UljkWOQ9L7qpojSlzWkhMLvJ7UuaP6hAt2xBMCeYw56NZuslC0eTvAML2G6p1eFaC
IKmFmTtlnwJHucrxfzlEOodg7SPvikjznPg1aVaA/M7BG8sAviPW1gJoKnDG5IuV0n7jVw3aaaf6
yQeqd+Grwdew5T4Qm6N7Ia/fMLqDS8lhodl2cfJiJaiYrorDqz3Bz62YO+jkll53tTuz+jK9WiFR
HLS38crYrGkLRtCtfiNt4DuuE32XEJXT7ph9uNvkUIlHRfKvsZ8C/ke5597y4MFUeQrDjUcnI3N9
xk+FP7gqFF1E88LcROIaJqybrME5lpURDmnO1bRvHimmbDa/9nZvEVpQmuBM9BtVvU9f1r44AozX
FjS84r1Jz49fgl00lUb1ndz5KIn5brgmrXdVFhTveLglzoixzQm57gbdNEu1Skc80nUFLa385qjz
/0FZk1ImtA/T9rTLn2r3hudXayJsgCVRQURJVz6NeuCoJmUGPe2yPZC7mV4oIw1jBKCpFN/lJyo9
T6BmVG5/nxnw7T/kcNszjFCk4BxW4wS8LNBn1l+uxyVqlBZjgRa/Myiof7Vg988WJt6w84KxJ6UI
2bqjsL+kT7oVr20VqvgTLXfxZcwhcLxzw+hnfWb28ncNjpT54tKT7Er+oXZDWy1+BmoJhXqmb79U
AxZ5rh1T3nJcLWa+ka7EPmkXywlfeqwpyXs9JlloI3NAdVjvzFNFHTVMuDId8HYu6U/VDnLynWoN
A1RJVaN/sMqluPRwRyZzhhY5S4y4sKBuHT7sVIwzOL5qVfKamgkQv694e5vrsz11am5LqckMrE8j
+f7AkjHomAUhYHhqBl6wtqQ8v6wAvfHmkQoGySaN+XwwPMhkgPSiu290ijxiZgtt590nz3NVRTC1
grukSkiz8tZXGZbzN/YGcFiHHOePx7z5myHNldXUYIDFZ3L3vtcpqqTWM8QK9A3XSsLA9hV4W5RH
gGjq+xGK0+nA4jc8mRwKdanbMNwVvr5BDNYjKGc/4xLX5EScOf/Rnu8+u9ij1g4oO82CyCGZ0a20
kVfPn1gCw64ITY54Sge0Y0KtOCbgb0m6v1poQny5/Nh8sO5ViWjpsHxn45LTiySOsUwkzALQ1JZY
jIBAm85I+3TqQRjgUg+5cg7gmIA3V0RnFM8K13/C0IDaG78SPrPcXDD/TqPS/bH7GSKlOSG4jzxr
eIsWR+yO+rs0aISeXRU0FAnoOdr5Qj+/QB8SgAPHWWf7ElZ6BaxdKStePFCiIKF5FEH8163/FoSr
fdCtlEKHI7rglQH8j2PJjNaBKD7Qn31i4mXtDgGfPMVvRW8QLeZraF1BSHfbiqn7AusJAcwGwONa
i8a6IpvGqvg/4jkudF1WiOwXuAeaYVNtwAoT+hCaFo3H9UNUF9VY8yGiDcaH1t6310GE9XY+Vbn0
hXaPHpXfN7+XGb0MFu1W5sjTangE3MmrCDiLmu36bqkgFIiXge+U0VePuBr0zq384dlM3XAgEkcc
6M6tl72dQkGNOmzcpJQ9M3mdTeo3vBLe7yaKQ545C4zsiK7AuwnxAehJUDYQdyolgvHMho7cjzHn
qjpntbWJd6DVWpT8fmARUy7xeuDDvlAHd55CSzUSdfm42lfSNBEUTTRwgclSwBisHuf9yO58dgjI
VGWM9mRuKk/LaLOnny4n1yuhUiDBz7C8GVj836WiREkpAF6zqhv20cM5igXPcCDowqOod3MyC/S1
4HjuBiP1xTbBdX7TW/cAJZwSWhN8vjhVGmUae+K9tPNns5R8u83Lox4goo9DGi/7ODyc8aq5qaKw
38D/Pwg5LAEtb8ltWMPyXfJNGNezQc+DUKLgzEdi+X0DS2ArJrkrdF7au58YAfnBg0WYIYIHZqhT
mQrEnLuP2QlVSavRC6yAPRywt/X/Kaagc+cU8Gmdi8NyN3XFKdauVWUwRyMfwnWoJN6QgKnEcGAC
mzPNEb8oWRcElPe22ihU5WOadaBU0ZjWoDk27FAJ1JV+WKi3eRogj8gPqlnOajyxNFXpAtVWHF5g
8F5LVwvooUJ8rb+7aQi120BUd7KyJOKcXzUX9rCl1Lgh1ECRueVFXdqxafobqBti7eNLfekptfMf
D6XMBonfWp4injT1fc1G4Pa0XEJOAixpsavHlKnhCBfnED0cMZ8R/GV8QWQB4Lzz3b/lo2MsBFGo
IN9eOFfvRtxTufvEejObbulS3IEzYT/Xx47zfWDHrMXxLHOkjNyYRxL2drCmKh+WidrsTAP7IK07
TIurjw1d+AgNE61wPttjgtmodEQkKmlfo+2oqIrDA0OC/1H7H8mIUI/FBSf3ThiQph1VE5VcvO45
/zE7wU0qBqpTdQgLnJoWz8bBL1BjfcAPfific8xRtdHiAycN+YM9fn0SyQAx5WOCABU9yJ6rZnO0
5XN1yxzcdENDZs40t5vlDO39M2cqYQFv+D1hzQHzZsa3XUeMikCwoj7yRNHBQ0PgY3FeInNFMdmn
oGjTn8a6F8uHrz6x8ymFvg8Ie+rTxoUplIZ0G/9HuyPlXmHN0dJEfKqYVbJJoUtvMM07gbe9SwlR
CorxkJVWCdkP7YJgRRhiGg/Sf/3zB7bunOaAr2KDSWlc8ndKwvNrQaQnEZ/Wit5Rk3jBRein+H5l
RQefd6c1G8j9KuG0NGzHqY2/a6+em6DgkHNYoa92/M/EA+VtTPItgVYqIiWTZ7rdkqHaGIuscFtl
Xu+4uS0PV8axBH/IIOkNHF99RDJNF+/RgfkrRZpxe3pfsJFxNqlZuAGbPZICX5FSsZkachnyTQKG
/sj1eYptjauj3dAdmMcXBTYdY7mjVeqvL7DZq2UmHMoerxhH6Ys4EHQUbPgEsbJG4qEadQKs/kJZ
SOvXo1ot++JkoJSTzxhSTpn/gBiUIK2owKleGQKCnya7w/CYeyCLZC9Dg+GPqF19Zyu9ghEZASmM
UvSRePvBq6ox1rq1iCO20AMSqFwnodM4GJqrf+bfjz6kEckQQ/i/VOSILqMfAptIP9R6IxsIbD8B
WPAkH5Au17jj9ZcVgygo7hCC5KH8GY7wCCRnVKzVbz/iZm7q7IMZP5S/5smH6Max6bWtVVzr83kF
qB3ZAAJUUnKIyDAY6Q1KDcZbbd91n1rJuUMEceFD3v0gpUo4cwdFNQ6L8wyyWN4xF5C6943hM0H0
MdDpDLbUqwZhAEQ2JnB0CTeaGQl9J1SA2YfcrJENMrxCaqAo2m1WSspdXuE+quD3Dszkao/vt4WF
7D8jF8etzuRUuQy0N/bChZv8qF5tYkfVpH48adlsnpxdBmRmkyTTM5LA2LrZnrsbcAPTh25fy/Lp
69kfWP3Y9jyr8DWBIfKjal13648V0sYTN6d5SnPOuw6CD5JD6uQD2uYhfM27PFU0l7YdDphMMBpL
T9xyx6jY5zmLDtBq3fWbE/+FM2dm0fY73/xvTe68iBG73/u3hKkHPzihCR6IyUevyTZCa2oN6qOB
h892efrJlSEOy2Cf25CNIEjEhYfOt27Na1cJJalczgNZksEF2Y+W5viLJ+byZOC+bXmlojCzJsl2
GG6zU+ZzX5gbQy86HH6zgNxeGP6PtyO0MPYaZeyLq+glTo78Wc/v6cEADLcdLE2fea/Cy46o+Sg3
a0oneZkcNsZfdRSlpod8HGTcoGcUZS6kGKbbik2P610NKx8//DQOMxSJPaNLyqw9PtJ0oqJCMKvN
NbOun307//nvg0paIqMgd+6EsS/9zm1swZ4chAGDx4b65UhpNEW3HZgwsnTA05LoPq4NtvUZncwr
UlOKxdj9iZljrfbgayL4S+L27RoB9QC0tXrZ3/pmZnLFKX5SouPKfGIPsQ/A4iqfGi7T7C9RAS0X
lTZg2A0i5eVb1U7QX5G6ZeoJfmWpltuOR7vxz8W+ffEUgsE+IzhXAlJJcsXi+bQlW08ia/MAOJGy
d8ooPIcN0ZUdboOqaXtGkZvUNcnwoFTbyvAWn0PZAUzNy0mjzp3IWGPNDPfgyn7J/Sa93GYilNw8
TbEix5bAMhFfVaVtF/DqnZ67W5vL+fhWJpZTk086O2oK6/qzmtPdeUAMad1vTlMcd8Gj6fAd9U5E
7SRAKL9dOmhAYSZJF2mC4ILSPf6VQhAwfQlCoYlABMXMYeAp75Cv5vz69mhjbOpuatTXTydyyeW1
NbFnnPTvsZ3xqtdPwmKNagJc6vqpnikFSJ742KrI005fZ7PpvEro3O1aoF/3ulf+//8mkTSMBZfh
XeN1/UOSk5l9+8BwJjW3YX0iI8ukBU6Vsj6aBij7rjU9X60QdRXVtfXST4VDYa7HMR5xjWGORNbB
v0iQckQi1IVJOjAtHuak1/aQJEZIgLpRe1ud3C2lAwmX5mypAyf8mD4QQkp22FU4+1tM5k79RBdP
g8q39s8Ka2Pv1sgFkxWCfcC5Aqjw97J94l9uxb+OFMcOtytrx/gVsAjaauZrVo/P/4kVTUs3TQPJ
GrU/1sKo8luUBJKPpJBuz6U/BuTEl8/sNj7GNRchOdyyHi1KYc0M7G60wIubeNeA6BRZD+9z69pi
ZgnLCx6aRnXHek13aO4ifnyI9MtoS9oc6ptFI3yE6KGO1tpL9Fhbgf0ZkjQ554zLV5AKM2vidqO6
4gAxsULuHWgZOQcZW07yo4fheoUfOTTOw6nUfWsbh98p1nNIOrzIIKASyZPdfuscnllQtFBPYjV+
z1cAO+b2NUSrIyXY8pnLFUzIBAucKroME8adgpmYu/FnfJZlZ2JftzU81jucaRQGbT5eSl8lfCOr
tPD6omCmPsEkO0A2efBZ6NdZDRZgCkdUnjUznDoFnqPNHmuSl5v0z2nE7iNDYz4xathmyuptOV5B
nsMLfHlKqFILobPv8QsIOcLHEx1gB7cBrz/OQQ8ns+6XY1Dfkn46gZGg+naUVuPpOeN5vNiPLtiA
8AF0Hkwe3Amf3prlOmCVAGXeeF/WvOSASmqVQrSHHZYPSCRhvw0INfKJOLaH0OeGVWyt3r5JybjZ
GfCA0edZMPm+7c56fcsR1Edjb1ifORw4O44pZvULLqOOONAfaXGWBpVA95535pUm+UxMFvWZsLxA
364pk/LsfeC/aDez/IsUFJ90c9029fH3mFMoLZs3dZfkrXzcjVy+Kbw0bzv6ezA3r0KShPZfcTHF
cCJRZxpJd+UMkGUEVRVfHCOUqhhznWBMxprSjWSqRrhzlkcsiOOQ5LmztN2fp0DaGgwejIoGRrZu
SdBkicPFdNdQmbFuWSAlg5Ceuq0meX3a5Q5lruD1u33sbN4jw9FNc3KKp8iZ1u8dLYe6C0RpLt/q
SYwU1CCYVrDzlF9qB8dTo/YWt1pV5Lq316Yi0MUSBDbOWsRuyUioiA8HYyUPAHZOB1OtZ7It/1jL
1bLczOKuGEDwPr7RxVgWvlfl7TP/4pBBWgQ1WLfxnwdGgNg0Yhf1Qt6Mv1uGMDJ7f6tYMEdUU/gH
or0lf/vxX1cbsb3Y/mnOQ/yerbslcGCA8wvPt7Sxhnej/H0Ew44LFVYO03OjNpepWQ9m4BwwJf0M
DdjI7JoYMxGlzDq9hr9nZmLK8lsMQoOUu4hynljzey0vJfCaAOxeJ/BXVV67Uk6T6UxV3qrFy41h
u13lLZlHfhYafnsRnpLkUJN6S4w7h5GSrFSDG+EzRtQpAQ8Q9bV4N4zYReGSO0v9Yj5otioifmLN
AwIIoRGCbDvDZFi0PGi+w+36qXe/yLPwf9lpHIwT29FBaPq5z9291i45D4Q/yHnTp9p+hAxlmqw7
/eP3qLzWg5tYc2Hc47mCYfLST5xWGCCbR4vnwmfpdwf648rvOq2Qv97UGvwkPD7JiSiEAmVLaxcB
ohVh9wrPOrRVO9IyqXRl91n0Lj5sjWq4pzs95bLD3DOSbo38YlGo9njut8xXzhw5KgMNT0+1E/sN
NjRP/MHzStHG0VGyvdmVDDqUeWxs/oZF/6vEXIlxjNFSADyu8qZwjFrYrCwna1Ua31pQaCVwTIyr
fTy0ff1ZnnZUtSnVpG5dEoOGCPTaTMsKN+x2a8C/1L2O39slKTrKfrVoBnqBTmKssJH0DwgZW4rR
qYBVpD7cjgcFMGLOj75mbcYxPDc+GEKFfCoFzlMNSnaB7awLQHhqNhBoAm08SXvj3sDDTLVnpG6Z
2Enkh5xqspuq9ayGjTST9RzNTntdtgzHVmVQVOdkFhcFzDh+CmkUgubB07XlWzft0/5hz6S2P592
69JBWX44427YKClpcj04eUvJYhh1jIbn45h1RLKJu8BGxPTRyv9KhZJblXAhnNFwMBmQzCmxjDk6
NcarAGb/xGr7xn1kA95oF18cRsC9nyxq4z6NwvS/4NNhfYuUHl53vAf9f6ikFS9f2iKUWLadV2SB
ZqBgaShc7tnLxg3d+F7uo9KV8oh0sY0Bl60zyR2+I8a4gE0rP653tWylmZvQZ/zWm7F5mS+wB64h
hDozt4zDJa0fvLd3IYzvWhrGFBsIqzz0mJLAlhifsj/l+n7bWB9TTaY0psjITT+eCFPD2jJ3Z73f
U8yKW7H9mCVJNHKrmU1gU5XgVrJI687eFI4O/3WPuQh+8SHGrs1Vge7YndAdfWEgLg/zWbTCrys+
WvPRZRzS7gg5CXsdWa2ED0gl3pz2SmZ4G/sBnECbJJWaxPE1+Gos6CXsbq8/IPAMoE3F5VrUbRln
IMApit4LxeBXghJ3SN1gl5/haUTgdgy2MxMDGkFAjnTFTrQzU2x4hx4BeQq4basMtgiij5VtBBsu
siEdiXTD2KXw/SBzR8Yrf4Jb7AoyTaQVeDiyJSgwUDDZYoyBkCfglW49J3rsz/tPymFrNLppFAme
T1g65+cEvPZ2Lfj8PvT6SF6LwJG9hhxJ9/xLK2AlnrInzF4h0TJzNrcEFIwJhZ/7Ix0aWRSgaFQe
5RCsrNfSnmEWqf+l66kNEyqHI1P1N4mVP8xcg3qFhxcc1OcAn5P7Kw5vAURF0pSZdEMW3407MWXT
epoX2dqJCTy/8CRX5cNqxtw1B3xhC4NaFM1Ym2MCklGzCHSCjrOECzxB5P+4+52FBC6LFKmKNP+D
VK1jYAZkXM1o1/LTrWU/Gyo3PV0VZvw6g3c+vu+w65kdnGU4Ke/z5ivWFwmclfa8q90fWFDSeQir
wvtgjuh5wANef7vNaw5xjyhxT+g3pcUxsgilzA1AglH22Scx0PD1V/+5cdOIYoHl/NzUxtDTkZ1d
0pxehY01a2tTfPqjf7hN6DpjDNjO0HNntydXEN+oOBB7PpjJVsyxOyGkZxz/NjxQKXwc4wmF29Te
4q1AGqyb2SWHbiB/y/LZbzOPJqAYO24FUCV/Q+k9YpQdhD3WxJeAjG5TBMBPJTmc2y/v5QfE7Ej6
GadNIg/kJSjBDl3VjxN7NCQp/Kfwf7h71sJWFmHMoyqj3jDoGeYRKYQnDbtIXoseczYQZrlbiECL
vaGGLwpmtXmufRlvRvbjqgsTisXxSV+6eh2WVl0oSIrPVIn1DN7IoM1lc++FBSoFRPv2oAsluHsa
7W6gmodrn9DTsl2V2/A54LO5vavCV5S4BRKrPpCj57UQWDZ06dJ0a4nOsk8YEOkKTHGFcAuruJbh
zXjChQ0Z0Ff2tsU8Ay93+Hs1lgpkwiXKFGVnRbfn3PScjMGCuhQ8bAD/yuScfLDWPWQulJ/WeWjn
LacVkVeNjzbaVWJHPHF1rOzvmF61J91+g1aJnISlUnDgwGzpaBVaF13UpxnoIACjwbqRzzc2j0hh
RvdazHKF/0nwtuDYhBFfiX6ccsvTwiB2mEi9mm+NX6ZoFnR/KRvmx64HwLd2OrqkyqbPcD9xVXLJ
gAwWAIkiX0mp8vlLKnEVd7GZWPoZ6nUj2x8yY5HTc2e0mNQxB1PKCkIk3Itc6tztNHn6SSNAJbNA
kd43l5AiJZYl3CM/rp5AR13GjXcY+fcjHddM3eyoxSskax0oRk/OfA5uJkgOh6+cqf9aaiK4zYPu
EyVLeqnUD7SRO2xDI1pX89OT5EXpyiKhMXKbYPIX04zlItRMo6qA/6dQhBhmK64o6qFEBPvJEIbf
qJ3lsTHX9mhSweo30vHG44QXFd4Pu5FPKjSsiN4be0YcZC/veLlny1KvE133AzPB3IzkVomcf9Qc
Wvi6d2ou7kdDtJZ0wSfgwRQ6s2/S3D5CQdvE+5QhY/Pt0HovgwEvfJ6p6amKJy5UAdMc9GJ5iygZ
tHFSGO1kb0fK57GTi6iGdxPgsy94132HRrlLhDMbfdyBhV92mnfkUYh3SDeWNgPGUKqQ+85FPZL3
RDh5ssxlSGf6MRBF41PEXshAYLGLjlEoaxq7oLeR1hQcCGBm3Rc9KvGfAaF9L2FbWBr9tyaC+wYd
6Et5l/CEw7CE46xrVp84w9TljacBLMupEvoTVIu5obUneXDHgvOmqLXVybk9JW11od94MCRIfXtG
jT9aAfxEtgOAP5fbMJDF9ATip0SwZdtaZtJFW9cdTPx6VoFn2OueIEUvZOGsotU1fMEUe/hWZNGa
cTbgTPnWRfrU0PREA6SG2XeBYI1erwR0alpdsPrcQP15NBUYXiIG9KSqjlDTCWcEplnSWfpHCLHr
ZcZ+IDNN1SWcYeaf9BardoRDqmjp8AxregbU53Hwwguf6o40k4VESPSzn59o0oPJoRMTO//z8U/b
2uH2lWEMF10hOQ9i/ZGlhRwZE9179FWDgI3xD4ig3I+axe6JmAbFI/nhKbK0bQn7idrb09VKsEID
UT4gB/t4TOMCghcplG7eS6qxUw7F42d1q9nfqhB7aZWTdjBG5BHN7eWak16bPyJyyCA4ueL7pXkL
Wdo3cRexAGWA9sQn+ekVTRvMOMFNTHnhzL43eP0Qbm/57W0OI5U9Cju/2WnSTzIgADUY97QPZY2f
sMpBHqkKipx0eXHjX/jFbDWalft/XC7Xx7hYvcB73OTb5yW8/c6YRYX5/HNrcJ4O/t28f+9Pe5UF
AmLJVfhKW+MBJG9qPMJIHWr9DuZ59SPBzOpIOjazhBafnKE0JrOBmtccpcPHX1QJwmQCnZLDuBXx
nL3+WCt3a14JI3twUNyMfO1ZGhwWtCX7XZINJl6ISfLTgTiPlc+o3HnntMtF/wlNrTEgD352Hbkg
otexXvVbuxtRa7GX85Y2rjITnybp9/TZLTL8nwyxxEnfJWsp3qkpb2mF3s32HJdrs4ioeJUgc941
iEYcByBwOvwPZFpp/xYt7AA9pu/UlTq3Etuyu5FpuCeP2sZzPpgjLXtiVzH5E/2cs96iJuOMpRkV
UaP5dl7Xtrm5F4dCq8nuLHiTWtfXxymPW2QW6/bWIENnMUdKbd+na1UEDIZ6P0dtnzQ6258f2k+k
MnIAvu3qS+Oa1vWQpUzYwkIH8mxrytLAsid1xVb1lB9KX6ZyU+UdRkkwf5VyD65QLFTvUhzm27Tq
tDGOwRbndqVeSA86Vrb1/7ifUO9W1ii1MSTeUqCurwCsttEs1pt1H/tZlnEWEzWnJdha+hD3tib4
45/IlnItTmKt9+/cGlYEMRzI7Lnne5/s3660++zdX2dRCvZP9+s+JP8c6D6hNMp6rvVFkY0GA09q
zbS6mJZ9ueuLUVA4ACXHhl4V2RIWoRx/3kPkJHQ31us3fSUb7NhE7bgZOFetoiXMRnTKWX4dAgHB
8PqqjT52GfH5JqDclf9Hv3b1BCbKRSZEmQnJEzPoKDHLQKtKTcSOAUMuREtMNS4/VMZTes/BFSnB
pGPuavI0/TgtSr6RPIf1QXyydIXP47il+rrMtecPp/PyGFeNPLCCDDUK7b1ICt24+QyHrTBXvv5K
YYDS3N8ZU8BAcP2f/nBmjdkW9CXdf9hYkduvXsyvLq2AyamxAXmWH/JsV4IpN/LxYzG4bENc7ybx
DkRAhnTu7scNwwfCYjGa0+XTt7R/oQY9KFaFBnY3REMMXhOGGI+mRuv2TncySmviNeeKzgMR+2h2
BLzX/woLp2QiggBagZxH12D+SWqyH4+lF6WrgOLmGchBPBlItI1i9469kt1SLGYW3SAD9wFjyzoR
oZy7TkDohfSppiwMRUh5ByUMJq0TBW9WTNwnJQBl5AWjLfrR+BLgAUqjNCWdswYBhNQE+UiIysTG
ymiYJcu+VBS0dSJpQP5QjSXYde9z+daM8eq7mrlUkDmwyu5qYHd1GYNd7ztXnyO3ts6014CNQjsW
1Wv0kU7oHVGO7HbiXrPaKfKyzYdXpVrPf5u8hTn6RU5JnX+oinesww47RKF5jJjoj3WwOqp8DQPm
qixslSCEkBMcxZpTedHA0+rDILhnihvuiEwmnNs9AieDNOqWKxeRuZz56oLdC2enf7tLsV2PcowN
BWi/pX+szzVJVRVo3b/4IE21gZcgxVVM+O6FTxLYOqxs5kr0Dab0PuI6KdKbk/ALyPDjtb8dc8nA
kpaWdsN68WkYdSJ7GbTkXu68zcCoBlqpcabU0nCk3RNlAVyqEHD1hHIFUKPCvuZzoNxTmDuztJYl
Cv3trV6VQzWMfiro6J3rpsOm7TohITOeozEwPSYsIcd3I69GiROfxg1iQrZD/wDDOwMDGkiyvuC+
2scv/2Nq/1s/bmsf15AkT1Z+g+k0symkp8jxVqzMLnlvPia0fKbaA4bLiLl+Pu1Uq5VQcQHhdDvD
37XYDq4jmEboEP9OiKbftoO+QqpO5YBqXP12qjWatLdsEnGRXpv66SeNLijODs+0UlYCtKuQ6Uq1
patv1XnToawEsWTLmPehFNRDE3Fndoo8kntBkcJHqyWU7mIUir8PuqIKKVnvCePUBhQNKFK9GEG0
eqf+3iJu2YJlE1EnXLpT+HDdPoLIeyoIxPr29o3QwYYIn21N22Lo91ljy0CAWxxA7D2dq5tPR7Ev
R/9LB/4k/9eOfycUgk2P+nThIIAGXGJKdXCApOxbOW2xVywuLJgmJhCXoIhTEa6wB3FbtBF6fLC6
E0zpmQ3GYpNoYFlyL2gj24nuywLw6mz7pf4fNRGTuk3jkarY4cXfMNo2SQ6n0U0FQZlBwbNaNFOa
RFmompsdC+Eq1heghxJOmEDk0M/I7Lb4EXTo/xmSC1yGPQ9H1sYRazHDe8XV1HmN2b/dOttPZfG5
dwexYvgLHsOYXa9UmYOumWauinsyl/Xy1hs26vQmDXZP5hLeq95T7qTLscLB2nZH4OvgUdWRTnys
5yX9UnfiJz+ITS/RGSB5RBcmhM38JNQenrh3nTvokTGZH4lmJAxDgOSSHULMiIjhusxV6sbhRdeu
2CmB1btVgAOrp7ishgKyE/Il1hiud9MhaYR6gONBYFqO85MxhHa4X5g3h50RMWafo4rrDuceeHaq
GYUbCe6QP684ssX7b/l6lnpzWO//SAkZO/Ra5auIqs3UNLtt1YZUFcAcbpi+KPCIUNCpJpKmiQ3P
a4UrcWQhga1i4fEyeRJgKrwb8KQBWdYg1hNXvg6tvCqUdkiemTV8JAiZIRJ1qnyqPopSQXR8PJP0
pNlOTy4uYNyblqH6PU4yzdziNcs8F6DMFnGEgBLbCc2XP4QmJ83sGNGNU5vu1vXtrUEBljq/SfDq
9Te8lDYuT9GBzRxWwK5LuNVaEEgdeXSPl074C5df81nM1D4F/G3qeDpr/iJt2zBrfPO2fOD2YC4Z
WOC19azQWHgFTGIWH2LVv+CDjTUth4mjCKzt1HYzoME4XQaxtDA8pFxW+rMfeWEUrsk2D9Ilguva
dCd7/wGR6RhlHZpWnTNyeBlLLrpIw8QNd7tsxRBrsHg8vXZCAzTlCyaIVZwaTCTMfwmbjjcRLvab
uRiKs4EzfYGZXwOj8a/o/kAhT/9NXJIzKvsFEnnlHq4D/jr3wk4vfONZrbaO2b46+c++VAMIYabx
5q5mdxXoPBAiivdmvAdWLvUQ/pSDVYl1TRt8t3dfyIhn/Q+Gc9pGn0Qj3L6nTo3PCvjUq5x078so
YA4/Gv82kl1Y/VM0Q2Doja9UdZQVtoKVy47nt3ZOTycvFdK9OLYo491rn246YMRTVSlFJfuRqJki
wzoIJvn/21TDHhHi2bNIEWI2nbl2lvkoYYdlP/zyeFGJIizVp551GNsTUwiMVYSxBwNvr/F/IUGJ
sSCt23GwzykK8YwodIfLcDkonj/4r/d90SYSlgALWOPXf4bhjfteZIilVYDfxjlXoaBkh1YH3k3I
Yf040/0mxZmBrsWPTdieNVusqdfsHhk1GqvHxAjLYbAu2tN/8NnMWRlQUhWpI5rh/k5McZtzR7Zh
JQBnzXF4IP2lDgra4DaOdtX07tkSEy+tF7tctMfqsz77m9ZZzV1IM/P8SUYYGLwaAYbmL7d6MYuw
/17ApsALM9jofTpafLr+IBh2FwD/ozs2YF8VTHSNsDiGCyYLoBokyBLFa/NlR3PJVNX6QQ6dViaW
2gZ3bFPY5DYOwyk5+isMCT3vHMIs/GbSaLSIEQDxPGL/TUAFf/0h0anCASmpOc1YeK22uTikH1rz
QY7wSldymkYVYX0vHPo9bnAOGkFL/MZz41P9am618d7wlgf2eC4exrkmBgYTOBedJwYVpjTxCZO/
83Il5v63Zk7jMsqvhwHePJKhNR16Xhx4zRe/rBE0WnEtapnZBSN49Ar1Xb5pomVPzRk1MiCI6Ssg
fQzZ/U+G8Ey7jW5KY5hK5DvIS0jCGvdvaK9GnnfPK3cCdn+w3Gcyje7H0DHnixW4kFtGuKBq/WMp
ypfRqevA2picURKG7TA8Rs+0Cjq/DxtZcfqkrfewA94REOZMGJtvU0+Ova5z9eL/HwUHRs/ASDpj
nZvMpa1EcEbCW8f+zYVQGTNZu4eqr3+Y233cQLnqScw6UmTPVaNQFWj5rK2ryOGhxbt36C+TICV4
OktYlyHfepVdiaY5vMAHVPQT8+O4NVKbd/CSBVmZgEQPDb4VxRCrZ/WRsLKdKC3zOhg0OnEDtrH2
wIfX6Qmd6uUMXBrdA/7AyvQLds9oHqjPzF97PLZqfrlmJlI6WNvU1PPkamteHPebIIjwiGoCjdX8
xNcgj5p4iOCahN4fnDk7Almf2FBd84Zeyh1GfXXjCgw3i1tygaTBf8gRBKzlWKZSAUhPaYUEINQF
wypkCElD2CaA6Svzl4fdfkKJc61bRRS8S1kpUtcGch0Jiw5RsXjE7HeB4wcr35VSRXqX9j8YvXUs
zD5SRbGLVuAoAwjvrlf8FPvo7R0hBrqzg6SWYGR35vOV8a5vkRQ3T3/nLpP50RR0MF6dkL/K4Byp
+E3qdaYlAi9OVdRpBt7JFoE99lgsTkALJsJihQ06hsJFs1zv3GSmXZcAkRtobuNeu8S77tpW+bqN
P9j4sBsy85BLlot3ZupnKudyg7/90X6synMJAbqC9V+1ig/qFqGyAXWcXwqIYveVFTFqheC1CGVD
zpI5tpsKr52G9iGf1ztd1+yP9BZeWqGrLPFJipsv5NStD47MbgQ3cbGrPvWzOrLk6bqkZJVST+hH
/mkaHxYqcT7Wtym7HujB7Mzk8KTA7f6CU8E/9NnFitAvVLgD+0VGGcEuw2STa5hrmgE12y+Q8m6Q
t1IEfGGkJXzMK1JDGZHG6UvbsCExC0DkYTQMjCkbJl+TJjnv5wgZseAS++iesFOJGojj38/kId40
13jO5VgCXSbMb73mp45lyLvZmnVwTZ+H85A5o3PUTqjzbbgIPyDHWiaHMAnT1dDrxSKhdFW0KG/j
OvxFkVOt1u8brdeKubMoEAoqEzDiraedibdz7FFS+fWTi7sedZkES+jeahL+Fzv4lu5Uu7ovoRYx
s+nofvKR0LVTbqdr9zX2Ll5tAteZ8wP7RCqxvCG/A0UzznaY8NqxuBsQ9a6z0uPlswvw96nsLZmK
GgWASpwlehJci12R1a9JhamTEQ2VLTA+6WBfU0vSeJjkDVbfjimdLJpxX1NLf1RTUvCAx/d3rRd0
5T29cj8nZGEESIs7TQc41PyF6Xaw0q2TYVV1iTIB3FECKwwzTgr8GKx/zSnMY0TvmUrMHwT+u3re
n0roPSadvcWLP9mTXAW/izrdAwZmK9b+Yh8Cn06TQHkTGHSMl9x8Detw9nqowe3LkTZ9jR0WxjMO
w11r382y2YMEWTqjbKHg/gJ4kmK7pA3c//ETEyTbhviPHt/jqhhvr26mbMGQR0Mo1CtGdT5Zvgv4
bhEP6NdUbI6Tgo6ui+QhKeQ5TlmJP+eucuSWrkhe4hLg9ZgH6jR5JqshqkkNZoqni0EW5WQ4yt6g
OvVl1QAAx8SAm0xLpef3J7vaFtJMhc7YrwYGO5wqEirxhaO5SGw6gNl9uqJ4a12LaewDGdedGGsT
mdTy3wG9nz0uWYVlDwQbZEWumZjwg8UTjibsO1w3BHydywAqRcXb2xu5At1/Yb0vxYUTVU3kK2ee
l0YRmrrvZNBppaIMPK/ukD2KB1y5EpvCo206jHL9Qh4HBsZvQ9JvMidK5zEbS944fIbapvL6Gzqb
C5HHihusIFu3X9EqCyRDvXJT4z4Y5/T/a/7/gSPuuybHd/eJS1p80Bbw1tTC0fGgHDIty7K0/+PC
OlsX2jnXLrGBpYP+OpdgGfPebPa+QR/Euvv/G8Ka154imSSjsIAEZn5JPSrDMP1JmJ0Pcl2Egqfc
h8WgHgT6Hunrguw+7TMjomYbxwFRFFA4mXcjDsgBspZqANjwYgH2mpnhrQXgyuLq3tydWSISTPfr
x3YkXfzvO64xQlfJ77V0u0qAFtkIlp2JrRQReMTUNfRBeXpKPr1VmnHLQb0+dLiDJ72w2pa0eK3a
1fPDlWEunmifb48uuXs+VvSSGrx+Wqdhyyha/aB9SwBJxwa6dzUHT4zfVe6KNj3PtrwX9KEwh4vI
ZmqGLxpVzKPhjAqHaT7d1bGetu8awRLg3woBIU1iqPqX3OdSLxkoxNQ0+DmtcoFx+ZC0eDDRscJ1
ZrSEJ9tJJnvnFKCe7U+QQw1PcoHySDWk0gJsDPx5n7miNmOX/wZ+268WD5n4j9Ueh7AHLc9aXNfx
NR80yi7+NybtolxL1GbVLwH1lthZkzql0guQmK7NPGHh+3yeZtseajkFAse/O5v/NVsuw3luo2PH
teSHjFpK09laKpue0qs0hvo8i4dIDRXwKz9a7qRts+EyL5V6cLBjJI2GFYQobMWHv3sVYMK81UOc
fDUE/xJS9qiPZjuAInC9p58yhVcOuaFq+jzHW/Ow2WgTFzXs3EffpOoxnXoKfGwxDZT9fBXImddz
RoNeIS37TUOdrqGXy+DfKIYcNInXN50OhOMI7RbPfzWy8MGSXL41Mk43Eu39qkEYBNLvT8o2Qa9c
dvLX5T9s44cKGguYvZUpT70UyhSdxyrVHShvmb7iQrC89Y7vbp21LuQQADlsjyjb57dmXboKHrXZ
640n16YmAIheBxOKdmcPFk2gGObMXfAsvMekXojAWb8Z3OIxlNad9NlhJqCBVM8gULZ1jGveFGyn
OHrVJSUvrO7l5R/H/E/7s9+KqIUbfA86N6sNLSuAzVov9RbqhdAvwkpLJLST8E6N5BwRPUjCAnLl
hrjiVecuUEBOspk5zVsAfFy+Iqmu7KW7BFBED2txVnr65ABgsW47kfzVdPaJ6aqc97Tmr9fRr3q0
JFqnkwS534WuX2VtgE3y9NJzQKjwNZZs+zNqkF+Nvx+NUwQn+TYaRWoDcvJvG1L1JxwyrHav4ryW
7EG1nXiWyMsc2ki2W+OZIdvlfntq8vXAKNswSyCTYSgLowuOtPQ+/QMbpZ6UWVh2HD3OtqC/uFp0
Kz8uVy4vwY9zr1xRNI78z7+ersNLSEioSamTiyuUHg6jSNt6IxhQssPsQiH5/B3JMdn3i/8CEz1r
MNgnd/OD06VynJYZk7hRcYt+jCFpnMdimGJMY6KEZg2DFWxoC4MU2D5yn/Jgo5n62v3YUZ5GIAPA
AQ2nCa+TVRtSzRC70QIha26dha4DF1WtrwOiR4u7AouCfTFCOVJl1VrHOEgA0yNxpPartyjWXEqe
N7eDOrObAUwvRu30w8XGPkYrnOIV5NlMDoXc3IJv282shtLPOZujM+WytekaxTJ9O24+zaoP02yA
e1tooqPqF6gm+AukqY71XSo6RJ2BdYp+ViZWmhP7rfsss62hJ6s/XT6N5srZxteN00vGzXx5Gw3J
c6JkJQ0WUarYKDRPkER74geRJ704UbsBbyBywd7yuwtv8x5yrpLNsUbdTOIJpVKfJsUvsxyYEL8f
+WNz6JTzz+zxDsEX1yVRH1y3mSl/JXjLw5CLkj6nsO/axy0qakHrKsoy0Bzqc+rF8faPHo2EBOCq
88On6OtKS2Tk0TchYhzk/21+eKlr0aatub02CET+9MfxTFeB+l0jgKaWnFDeX11IgZtrydTshZRP
bELOT6qqBQpSqW+p/JRHayTmoGFl8/fU+C2yvFVwdXcYqGsZnTVj5e2AoceoGavp9bUr81gQdG09
BSyOQl/lRZxjc5XFiGes6ankgKJdoWmZW6nt2ZieHjeRMmE93ueGtdLH0OmfNpI2tUsQfXRbeLSk
Mjx0dvQDLYvAVlClD6hqQ8SyvejHxog113eQVPaaWO4RR4eErnwFGmUJcXzO8DZiD0fdNjC4W82A
/SHtmI7zQr25qdMPq50iVMqNK7Bh+BdbKDGCmly/2brygvWm0BTe7OPjB462wJVv9Jnhr4weWA0m
n5Fc0CUAQPPQ3rAuP69kiXcESD0/CpILFWN8oRnnQHzgGdam1F6mBaR54ovm60EUg26xGxqgAH6h
oyRLoRzasmJ+EZUkWvWQQicSiwK6H6meKjq4ssvPzsTqRCOiG7iKYm1W/GKmDvOd/tRmV58mwxXP
N4VboYkQzzAhKlqKu2L1o2Iz6LNg2l5oYAUHgIZBEjOMdGYnFzgzSnJrtp5JKbglR06/E+ksXcLg
CNQM4rjS2WaincR9BPx8Wf/0KSs3xnvaVGCk05IDDct5mdJuaVt4dYMj+1yuIxK3G86IfpORkiPu
NGS+JfUQ2QKpE8LOKpAD0nWI+T7ypvkXyPz4zS3TiPHcjZrNgpJDqvRhOgPkO4qDThtODMxd9llU
iimJ0wmms73TNeifkF6FoQi6O/2UIxoM53HciL26B4dOtMlq3kU9NXMZcZ+Oj+nqiPbbZ2ITxyXY
R9SwdaTB0Y+LSHUd7SXCARRCBi62NLftU/n3bkk7VeBshZssMenR1cELR8cc1KUr0phcvKfEJwpH
iaZt/fPHRv4J1wjLiiuXsB06JEQhIKrdlWOfhMYLSoPjzUa08WhTERUclbOQvLly28bpVGbmgPp6
3CMO0ampilOR/4j1zJlJUpybElNpBADO9gXH3j7HlJ4vJpRFvbvGyCKyt3IgBUKsL1U5bJ6278cY
yUiORuyd4a6UNxaeBxyG3oRtgYmADViWTQ1PQJJq5gHYG9v8qJOzD/L4wzMNAZ49Cw0AvVRyvpyG
WJZKrq/4U1Nrehtax/Rvw0dCxH6Ns1L+ikXFbXzQS8wchPayRqRIb3Wm/f9qAjAPd8Oq1neDym/3
GH/phyBpyOaeK8khga2enYSfxwyiMFHw/qCMuIc+A8TFzA2Fv/p+WNroJ7kMATssXqoxB1Bvnfz0
tWFcKmTLeLMRTl/eSPU1L6I1NUJJeMRbJ5J46RiFbsI9h7Dl9uBBBvMMXxMXktoFvd7hmCEMXNvC
skegWFwCsKNsxqB4SnmD0FzsRIRgEuvgxGVk/NnEX2uBwltQBv+ecPq37pW8Gc2rZNFKW5soKzxH
9Cbeupm7rundGynlpce6r/zbymNEBy8LzFQ5fS+tEkKzekhO1JLzprqNN+JFBB0qF3XdZdEuwBqi
5hSANwGorWmXnijEUw0haj49VoHDJCCBja1l0v+F+3ivYHi3ogwC/V7ZOTKYgkbTV2kzI6KsLA0l
sk3PFvWMA/4LsoKH+Nuja5/qeu0zDTzomT3nO9suIlPBHnaLkg+jMj6JYq6U2u2YiJdcwxAwHCGm
jmY2jO3wrMkhnsst/8IlBcSv/5xaesBliG8atmFyNMJKfPObjUwlixhQmSg00UF+WNpWCJO9l2XM
T9C8YUXfy7jnnegsLTtuYzzDYNUb2ndpka5Wv2StkBhYKnyj/A/KVKrrOP0iDG9FFpXDJNga+dgE
3Hw8oKeFxZzifNwirYqMXFYY2hvBiKYZsTIKfFGEz8Mt4nQYjhbdwGMWl8O1bEEjphpGoEZCbcP7
bSQ6+gTOZpEWYqaoqwbvj/GYcFLPOSb9QN/WJX6Jf9GjQBoAJsUeCYWBK+OGGbmg3uByAcwsarU9
lxloO3WOz5ORAA55F8Wntt9IgiHurtov3cXHlkzrxcfvFLZy4VsNHlJR2beJFdpey9RjBDbyM+BX
j9RRbGLq/hwHfLVZpFtycSlnIH/1JW85YdAeRH1vuCJBOCTjl9hnE4hn+v+s+IJJBIOEuOc0YTvo
Nd2BUnXEYe4C1prQnP8ZGvKSwTpPu9s13FFiOByTlnra0J2TrV9tN3g0WiUJJNx9OtMqvfLMXmDb
LySxutW1MK8djYkYY1WYAZyZZaZt2P7gCfJ6E90/Zv1cWH8Z+kPIYk/mQqMPLL10H3DlZ8NEXAkW
y23CE+hb34Bm0PUtBFMAM+z0d7rTUZURB+s7a776ETAeX7s2BSfVDGTDMIP8Sh77zDW+PfPQJRRb
h0bBOttdxqByvn0qF6hgzdI0+UePrT1hlL1ECGCHZjp22V+N8bA8mP2PdRkVoaJtnoj4qNDdcftI
TdR4sS/b9B753T4wTNrf456x3ip0RhW3Jd2/w0jH3KLtavrjJ/IX6BfJMQcDeS5yZ4BYe5iCEnBN
rQ3ioT1RON4IzmDf5FWUfdMDnsGLdtpd1wEQ3QuWyCzCJOdSZT2jtBCvFYAxE13nYSUhLviqf3ul
u2NmxMKUCY6FyyjKH0mQoddKSGSNF6+snKXp75iEWIgMe0Pmm+kOzYcyciwvWzt9mtaedX42MncX
wgNwJKUFlVcyMz01ySacbfkF0wO3D7Y69UVPhjQ+dyfXwLuA9LnkRfgCCf6grO2IAkOPcgXREtzI
ftpvdFDOZlnW7TcKWpOUFg/R/1FUbwA06lcwusObk9pDMijKxMvKCu6UNKXUhPJfYH+oTk9AtNe7
jNEj6YBZgxhmSlUrMGYT2BkoCwkDIUmmoW9Zmdndw7WU3CDl3trvxH+ygH1LPOYR/guXUrjvoXPZ
F0VPQpo4Nr0PtioqJSDUo0ICCfF84BAYkGycnmSRXvfFw+sswssQGQizWBdg8KUmB/psQE2yMSjh
tFRZaJBRlx6ro4GGLaLgIWcjvTP1MFV/R3RjqJVSh3ktd6k1gGoj0jfAy6Ll/L+JmMY8W1hhWJw/
QxnaQfLECsWPLBKfvPA5LfM2o11R2iWQIleg6Z9OkrMiTs1PS6YymOIJPPj97tJBZXt59QAuSh0O
pZQqxDW77kZxQHuy+nddQNA7sy3vl8K0TTt5zP8eNmIr6i7EZNNEoyEz+i4XkuscH0jIRlpCXKPO
oUoYqY/ydnZThAzc9WG8l8AU4AaFJkVX7HqhdoU0zFJyTtQkXJRvQ1im9GND3vu/JQOH7MbsVUwd
iZWgcKHZK4s3Gu8t/xnOiBMSh2ccHNmEWk8P45OVWhe1nJT2yiu4gDMOoKcU9PVVNF86d2jrMHPa
r9ZKd+XzaEFYRx+Jatv5ODykiK/39Qb+rjR+gYDO4M4epn6Te9B37jzfVGvcI1jMztxlKY1fr4PR
CDatNjKSuhiuNCnq9BhSxexGyHSdjCiwogq/C9yVqdu/ieqh0Q2TSRNq/EIuS0ta55sB0cQwQTCc
9vAz6brVzEc91nPkTtcj60nd0yBnuvqrDAjf+ngclNtuPG5MgcjwJjYDfUtqVgIfBi1XwD5vZvdJ
VhvQCno/ZvCN/HnmWpKci/7kCYoLx/C/dvaI/3lyngaleLXiAkOSEaIvFG0Vg1FM6H6kQaQGxlWa
PUth6f7BLhKx7OJAwPo2hH7Nodmn1peCo00ldJdP7nXvOzkqizuw9J7iOeJugzQ+fUa2w0v5QbrI
bTtSku9GQISpvdXELiEOFJjjVwy36UpR0kt9UlzjBNj9BBBKHQmlx9uNNFPDENy3PpkuuzPD0t0F
9qXo98GqwzqpFXhICjz3Rk6VU7coqqYFi3WZv6Ux5Qgpw3qgqkT97fZ0cvOwqaqSdHCpwO+a2qRw
wBiu6GrOAkJoPRkCXKHTEC6aHxienovSC9M9PJfOC0D2V3LAERO6owmcHbY4PXNe/QfRCpJJ7tyO
m+oJAmj18A/b3rm62fAkpix1dvIuCzoXYP6jAe4HHPmuSvtJ2MZCtx0ILNPXde6KN9fnrRop1kOk
7qglODyxYf34iL55+hM/Ukmp8vwhbbSJI1YaaF5/WXwSA7p4sL1EnKBEY6igx7SD7OiVtVWLuDIa
DNNRclEyE3uKEDsU+35u1s+Ku4VZg5qZQygQNpAE8X8dM7yzxvYj1TmjSN2jqK7JKQ+yiJwfZoMA
ld3WDaJw0AY3NqycpGW3ijxR4A2faHIlf1inmTjnUex+r+no8MGP5y0MsXRXuuQmHgJwcxwqVZ89
RBXVgY7pj1sJifQ8Tm95LzfyoGNtCxtAUf4O717m9ip9uUvg4uA/sPWldauD6Fkbxr4YUkXa3HSs
t2hs8SAgXpyWM8tWSh5onTq0So76iS2+XRMpBwg0DkYwc3CPcVOrQqV2S7c3leZIEZ9yzCOgVo9P
I+9u6Y4q11kdkyDZRX+3PT9kjUTvoteuYxpdaa/YIjkaRhzVFlqth0N3a2ojkNda3qcGVTyZiFP9
3493Sw1WV+1UtZ4mSffBTEyw/F8/sakGyb1847vP+kBjicNqde8Lpj6bb4b85CfKs13s5N4SPgxw
7BNuDhAyXomU67iySvUlPC7lUAyzj9kpYU2Y+v01B5Sj0E6U+pVDAMUghRdNFIqbaEun61WRz6Z+
7fAcKfaOxlHKZrQGhhKeToFKIGbwgwuxYTZHAdiHQN9413aaYS4GhYvrFiP7JF2wU7v3mEYjJ+iG
59OkqI3MWC58ojpan7m006jeuZVQ3pfbVTQz5w8JQ+6kP0c96V8bE7gDX56bq4XISzHrIRNeo7Or
fEpyHnkDa+ik7BlgtixJNT2kmxiBXP9t5SKtc+vLzcbjx4DZT3Y8Nft+D4roEh4GYNKbyLFWNpNe
8IHYplULz6jQ5PFVCs0jEk13YYy780+4+W+KBrutdyYZ53gygfQGHNsyWupU55N5xodUT7bX3+5I
FZwHdZwVSWsZKy6PAUOj6tsv5cytQHeDHM5Gn0u/dQI2jIk/QvBZpWLT5e813O5BAyBibz75qSAh
x7ySwYMaTnvetGEFFK/3V87MHEx97CC807rnSrM58GM6ahvTvLNfLzt56o7l9YZtX800TtDp7zqm
ZAxzf9Pt0NEq01yQHmNvw8cSocHJAhI5zY/o211RARdticc+9/Dm93z9lWikwPNbnJ8U0TottKyZ
HkhvmewpzwUN0cuavp5bcziQVsGc+1rdc37j1SD1kbu1yBCqyE59i/ZL3A0vuCFIXUbnaxNFwOlt
MiDcKEeA5GOM2Ivpfd/aE5nCY5C/x0LHwVpamoY3RC+TsgGYcD3fQlIGrjcwifZjLQHyPIemsrMf
oMwd/S4QYVldlh7IWgc6aLJSf1ok7y3eWM06E+OPPKGNsnIeB3HtqJLd/ZeXSB5NzInpdxh0yvce
FLhp0fIUv4/J34bpRpT8o80esxOzuv73PsP8ZHejkGNQffWfiUF06qWCdCv3gvYFfAxWRYMM6UXc
ET/xSospfIjTB/ck2zEgklpqt6wBClaZKEpmpg+enIxDNn03xoNtLSJyLPB68NFxiEGgYvsfdhlw
2JTlNUuQecmPHErJKfYkk4NIHg5+JcFrmkrlINmIhgtlZSGmwdCAqkCb1gp77/05uB0ZvPUC2GIY
fVpzjAequu1NMoU4dPfJ+NaRWvj23tg69cSrL3YKxLUz5Ynn0zJBt7VYgiJRah6Wtr7NJ2fhJKPz
3X7vSXH40IZQiUdoicd5Ht2ItAq9OZ2cIY4FrErzld9rtkmOjAvEgvkVif6kXW1NGAgsfQyQwV52
qVSYyoeV+uw2w8py5wNOutYz+UDfOSeB1QOvIS+wBQanyu4YlQvsQhPCiSoqd9DXY1eg5fkViwev
sLCqUx3sGRBEqZFy7BkkleFyX0HF3jv8G7VrFPxiRwVYcunvzHL6vi3NUsKd59PUrJb6JQU0rfds
fZ+uH5SeMt3slyTYLWBT5oZSlMi/wopaOGBEE8xBm2oxTFzczcJsQlFrm+Y11eWN+8y3dBBG8hTR
CtnyF52fN3HbhXqgg2maKftgNJzYnNwr9X1pEjdcb/EN5drgP49/T0rwhCuMltVEygGXYC6emi8B
3J6kvrZsteGN2jh7/RE6O52s2mhE6ATxImqvhry3qLhOk+iP8wwtARRJ+zRDRcEGOBlTjgcPTDtL
sdUaDNkeUK/N1Co0pRRKorsK+E5Gm10jzFZAERqUjvm8noctkApa73ldV7fVaRXxfklmfTVTJA9h
mcSuKYpvnAhnnR7U4Hdc8Vmof4rqrFeEl4hBgAzctc//CSsgpj7VXb7zwbhAWZLIbkslkytXWgxz
TbfgiNrSRU44/BuFE1nRgd3TBmie233AVt3QOP/WNTivCe6byHfSbPpeNUbG/486BfgB4Ioo4l7x
5fGsQC8gKyn9p4SfinHbZyj7htMkidu2k8cJq5dd9nBGENKg7600uSI5Zhkkru0B0rNh0Nr3akSp
Ksf+OUa61+jhyemtaxlKwJiJkMoymDQ5fYjMAaDJLU1klekPY6MTMrK40ytei1RA9p0NrMbOdYTC
So13r+rXiVlQv8qFeJq8fExB2D1ahx0uDz9iniOedmAC+7MaTA7oBiNFckYnvraKw5/C+hDM7i7+
uPFuS5BDKnA7sl6fQ5fvq67BkxWXrqiAk0I+H55V/8ZBZWoHrIpAd9m0OgKyxF58por2FOjwZROv
gaaPwc7y+EuTIKShB/HZWyRAM40arzHGQ+NB0AuVC8kATuhgy9FI0NV2fsZQhodpL2a3ONS6iHii
pjSPeKa1QUR7CV5rTUKCP8zvh/RTjdmKnkhrP3jzpzU/ndML6T5V6f/VW+/AvoXXyS4HCZsLP8Y+
sfL2LKGO//ocKWs+juGFGL7P1qmlFDuA44743WFP90fdgpshGLNQRcRa5ayA9SqdUP5sjjMrUOdJ
2SM8JczO2wvqzaMKwZWOvPFGU/o3mH8LpjTsLRb4fFd74WAiWyhyYq9zQ3M7MmbrN48FCJX4ZgSJ
RDjA/IWglBGsvdlB7lA5I2m/z5Pa9f7Y1/6GCH08BU01mNUuAIoluVhqEFeb/sZEE2UosdkFg+cr
gDkTDTIhgBmLpdGIEkdQAM/8sMxEPjCNxzhOizG6DIgxYv+1HRCZvqYfgJ9G5PmkkQSbpGKzaQ65
seuy9oV/bmS2+RUEzs1A/+Obo4fYSLcG8Qa7ObZQ6eXDLIaOBQQYD29fxottwzKLY6gzq+NO4kbo
CKIOUEntNHQXJVfjf6Vr+30odET5ULnDaloE6yj3uXTf3CSZJtr77L531aUIqIE6bnIXvOVReIOL
viWmT8U1ruzZimGXSXbWTC1AXR2ycbhj5wK6SB1jeRZt7dGNVJOv+WwDoOsiDRSkJgpj08z7+1rc
+9C1dpBzpyOuPJai5wsH9Qs1Qk80AfxeFRxvtA3z4VlNwYBDpT1cMBVXE6ibPfr5/Nx2ZwzNCP0Q
LHv+3CZbl1mzJNrH7LeWMaqz89WvqNi80NyK93MRx+x2gARKmCxTqtM6/vAG3fh/kaI5batWpf0C
Wc1NiYYGTD54S7FJwRCAuBuZ08ONijn0n8/wgaNaqyxJ4AMqSXoZEZmp4DtR6NyQsiYweMBWCasb
ffUVdSaOoCPDwcZMJS9Aou5D3vpsGOyYkgvmxQuTdWGIA1GqvuA+LIxm/Dr1ufTzlrZbRx5v8uJ8
8Ak99p76Zh4COZznMswsOsWbztfGI88x/tGQCuSivLI/ACcS3c4LMZ2OJ9e6YOQq2rNSy5B+zDT+
hFL3fYBN+od9P8p8lb/8rb85A+LQkxDYy/8bH/J4A58t7sIar3+bH0fasw0H0sCt2XkkvzuRtr9w
a4LKujKFJTbP46tN2Rj6ot76BFX9q4xe53qnBC33obzhQQdqteKei/nYbAEHdmhX1kbvVIo3umX2
lEcEVbG+RkvkQm9B4yQPYoj8gWPRXLQSyVjaCSVLeaiVb/vsl9IO+3o2RZ0Hlg5s8g9Nsa6X4n63
0eYkmKWKap3wMcsPvRhLAUvEx0FbPpZmeL97i2bdRjes+62SUDIf/Y1msbFh0agPMLteOYS4iAwN
9txR0OM2qNpEdxEADF0KMeBFWoqric46I6ID/Fu5y53Zp2SUl7WoZGp7BvEOMs7I2KOL8v39tLpo
pn+xLfKRg5rpGpC6bA9rDIqM9u16PArjmXcTcIf/TwUBpcpoL7g12kQctIVvS+xymABeeEWlHnH3
c+vAQ+5qOI8UVhx2js9gTj22ydiAbBWI19wsGxVisk7Q7KpmO+wmCD+LAgoOVyfVThaKsX147p2g
oxLUWlYdhLlQnjm9mRFs1OFS9qhway17C+O7elGVDrcGxM/bwyKQ3VPBUS9oIh+F5oNxOagfzqvk
1Nuf9blUOBsdoeyPY2dVgSiS/Bp+MVa53gC8K/ZZnHeUrX3hq8IYr7decfLFEb5aXpCp5LbcB+TN
Cqe7bSCSqbAjFFymRLkkBpH7g9HCxm8KJr484BMVSSzQJ/Xwn0S4wPlGwanxS7WIbRJlbNyomjeJ
RdVJ4jDdnrxgrhDWTSVmfiRNF43NYwNBTOklrNIhb7+euSiMmUkMbSrQHsKzl4T5T2EXQc7uRSTh
fyAHD9VJZf2j6K5XGS/ktekNxvocddQzMfyVPw7eR1dB+uR2oSJXho9xkWwZLRvTalJaF4c3KGLq
CqXuhInrS5RThZUxTbe2IAJsgvnYNjrLGQoETD0n8qNqj8JEgl2xFmtQ08Soe30EY71yb14Ecx0e
99tARi4YFwBLv7yUdDXlbpmHe+tt90UNWV6wuMP23FowH+fNfbEXxrqGrTPxf5hBZGKkk6E95Llw
xhmt6QSk5+k1kka8izM0bG94nW/0HC0Mafv6NAy65On+dN8rnZnPmT74uWsDis1OsjrxkWYOcA2k
I8EbXGdyTnxt+MWSdfmLslaRZxFHDV8vN9EbvRxH5fQJLAB0IyX9Av3eYptSf4837fYB66YZnuPO
2jklK+vMcMfFI2oyIBtiBCqS+hpyII/M8Bos5sd7tQXjqXpOIUIwV2mdBzeuCrc9pwO98yvUy6nE
lwF/N66+6CtVfTmh4MZxu4TyBxNYH1Tlu3byZWHc0gE3Jl5DrWmoG6gVi7QfOhonTlCl0uMSlQ4Z
yUxKoUjrWk2RvNmroS9cRmnPAmTViwZmb9QRzs64/6E3Qt0zqZA98Xf5NaOdufeFygoV5zc7OXb0
EOpWnxNd3hhYI3YH2awXX7ruOnUtOB2yKwXbULNT9idvpjfeK6EbetgihquWjkCTWiyQl3nIWSgK
xsb8dIBo4CUxufjyl+HYD3tQu629RLn2FN97YaLlxJDDdmTfIvEANVwkeDYJ7Z2nZD+7jxTAdFa7
Mu2pRBamdj1vpQ0v4aOG+fGIkYgwS98xZ5Za52oLKiugyrYxNSr6GUMtdA4sr9k5XiYkdvCGGOtt
8+gu28PQR7F9ZpvkVoGfQnbgJAGnnSCbG9bH2uzqYFsktkwvctRqeY6qBmxk4pzoDhoZ/2SxzAAD
wJtthhMd07D4w+13Uyx4xIhU5c217e18MXuNrIDIPOwvOwDpJYv2B8SOSmR4RxOOitGQVPaANluT
wgFI4pWhbF/j4G4EqRlaz3Qrfo4W8t4SAGf9Y7yb74rrCg9o/v3wnueU35Puqm9FVw9Ypfx1YKde
5N8dAAmpsWQ7f9pMUxKqK6CTbjIUXHw9Xfykf3+ydK7LEfX+x3Vdv0i5RJVwEu9TnKnoXQKYSgN6
LGUdaEMObWocL/yY4SgldNUBkuKjmRGlpOPnYn31cFD26/QgUl4IjLYPXmnaVf072RInUfJYfGOo
5FGrCX++HfNqBPYCkKxu6pgt9z2gyVSSZhDFMHHpX/VE+NF0wFrqGqc+9rIzF5tKTud5wdbRfMCN
KAy9f7hfvz5V5dtACRivPvRK9+joOcfzschK/38pDWFLfzRoCPruu2nqTQOc6seivbt14fDXbHOl
q8BPFDspKmIv90JM6wYa7gIfcE/gp0kfokciy/UA4yo5zuF/D95S1auaLvY7hOIrtczbiwULCDxH
Xkdu90DTFOrgw1NkoK98GZWOkNLDdy6GgX7cdg7mju7phqszpfz2eTVAjT9pvxdJPpT02sedazI8
PhSgkWbtq6kAawMcS3SBF6pNiYhP/WLVxBUYZgRj/FvnRrQjCwLjPXGQKfju9mb8+Di8yy+V+FrQ
dDoHmviEpQ4thqTHvqbRvJsA9PbJ+yA6iKtvsUWtYZaOeVc9ymdELdZ0Ts+Y2ioWUka1V0d5oZp7
RBIwcruaiquWbhOQU3eFfdWhYgQS1UvwC5aYAsL9wbhs2Y0XQU3w0hDEaWdv0kiCidD8Bz0T+tod
/sufgalPr33lKwHpsvJZdfWETwzMTbU3ZWhpYT/yC958qr75nP4cW/vDlKw5qTUqGFUyIfyHthip
HajidQe2MrEfYK01FtwF1etqWM/bvDiatu0XOCs9rmiLdGeRO5Xc1/Nz08cDBdLC0e9a7z30qipC
rmWCznYLzF/L7XaoSeSw2T9IQUEZ8N002F046Tlebl+85JjbhedczTfZyVnFrHm4Weaj7erKH6vc
EDP+oG0k8orGWEZvtOL/qrtxc1WdedZj3/8oLyn6FOPYbeEBDK16sv2iPoEFDqtYuUNCc7Zwmq4/
rSLX/a0P7YB7K+g+n7KTv/ddmgojfiXP1msmQAsdDCuwcwsatKrzoBgziPB7llA71kZdNa4/ZV8y
UCOKN6bPcayHHDnY/R6IJxy+Q/oUfALFc7gzXmbRd1Bnd6Io9P6APOAvTA9o93lT1+1PyGUpCn/N
Xk8ARoyIw0pKxqGU9zJuwy0sone0sZvGD+c0Nd6HKxpZoSJKf+JSHQNo+wfr5/S4Iyie76MRsfJK
wv9R1tgr31Z29owmEoScYVpRzoL1LBhHwwhwDlrqX4W6bfuJdSHrOmcl3IyWqTnxzclvFLnnpFWU
B/7fJryCz17iFPK9L9M6Nbc1HGh9YsGE3nSAs6ueFJdjkNxMGAcI0lmXXPhfuuRFwyt/sjHVHFVU
t9HVQOXTon7xSl70FoPbpN+sP9pLRCohFEemClKBA7NfRwBjOCtP+cC8u35j3YkHWJ95csg0HM6R
bWzHCNM2DMYDIIY4eJHPUjTWK7gjKkP+s7XD+NZQ5futErizTgNcSaFyoJa2QKZyRx+bVrpHPGgw
9Ep7/V8PhUbUhHkVNLt8pbXNdlDxEMDJOvNOLQRPsqKbzdJVLUkJg87v6e2XAnvi/N43a/WgtNo5
Mp71slI1vQP7DyMm3lRVo+43hJWcbhdzbWm/S5dDsvOq/PjMl4gRke4mzuPKr3av1C5RuccSg+M9
Grci9/IUfEjv0DQOIO+OAdTe2yrG1QhGxwUEfoLNRR7SsL7agDqt7JnzJ64HA2ZkGqsTmxEe1fz0
XOkoPd+6HC3xGmZdaoxl1sIXtws4ll64kFfRZIY/Rv/TzYQdgkG1vPGDm+Iuo65CWd0Wq74+EKhM
evEfoTs1DPHE95502EQKZePpmfwsGjEK0M7oL0uaiXZFhusTmFjMiyfrhJlAgj7Xx7aC90mUVPT4
qum7WFTl/g9B88B3/XPBPgKInripC5hcZeEZiRNZwkm8o5XL0wFDCHUjuo/ZAqP+ufdavnZhsx44
3Z5/Xh0sKAh/au79RS/DDEukjazdoG2aFn5VSYxyxZ4DqyefNXs8DOrmSa+fHuy9jcLM2/yv/isM
mAb2Lq7e+hO5kjh/NMMqXYxwlmLXD3qvctM+uVguDDWJ/lUFuWRLfn3A19T+25nk3Y9FJA9A+hAv
n05UCl76fHT+pi2fVS7mdxbL/o0lnkhlFgG4a83z95FyZxXHBRN76hA6PRUPzDawGo1fASWKdEi4
a5VxmpqKKJSH8orHTrdMEq6Uh6/WvgN4r+iZoaCao7sFnl/ea2HB8BdkVgyrkwppP1au3KjmNBSC
c5yhjIW6XA5fU3pt7Xo/a0sMv65Yk9eVi4a6H2G3xOLKa8KzhVPwdHfcz1OwidkoYckvpAb67ho2
l32L/ZbVqGY1zgwxmYz9zB5kfTu6ngypqtlIgj7aoQ0OykrsWrkLESXLfn2CcR20wjzRb8nffzuH
5P8fjNCz5fAhASuyyGjVNjvdk8eWgOXOOt3M1e1nDz5KX8ubthuS6Os0GIcXqI0tQbt1pSHIfUwO
/3zsJBEnUfZhV17b6nl73faAg0laU43WrLsD3LJFWLfn468tPkLhl4hSCThCW+qS8PgDnjEnhsPT
dP/+ds5ZxUuF2uenI+W1cLOFFLwmFTGSB6SYsvGPV0qvbofqaXtLlfxEc+lM22iArrOwwQ3M272u
Pb8bIzbB7q4mB8fW5Lacn86PcipXqAmgiBhZsczR1nktBeoO4ivAxHUSXwTYP03FY94eOU7G5Jq6
H0Ii+pGLTOWmInT5Qwqv5uas37ZJJ2ygRdN2Cignkb82MZB5+Uce1xbEu8NEF9YclddHugOyWMKE
fCYdd4JTDY12FS9T4a5XVEDQ9kUiBAUW6kPAJ18yQm2t0XqIj7xjhl13vE6wVlGd4c0a35ikTbtc
+AAC7PcVsvSVhVpeUNAAYstlLcjiTpeHR7eKyxDLTdWd5k0c6kdQLIY8kKe1IpRtyfINFoIKTPeo
qyaRvd+ZcsTHFCRi0K5gKFuoDm9oopS9sviF+XoGLb/Zc4+Wag7VQA+H3QQXteOr3dQbTeVOnOBK
dLW4EGa9tf6SSF6+4OYQZVe+8PPr8C7a4D8I5M1yK2tYBxGdWg52+Cr7VcZ8q1ASM5loGDCP8DYu
O2RLNY+FuHgi0uPJRK0jmTXErGho+k1B8C4hKh5d1Vtm4STGcxJth3EnL89eL1LSYXlmIPf+Wlth
x2EVGVoey0KDCsoKt5o29TP11xSQnPsZM6mUvYrA7tcylXBbe1/IPeLgvscqwuBY5SyJ3tlMEXyc
hpcpUkW+YBupdkvM2Ik41JyFRD4CWyr5EBXSfVOJkV0JspdUOylr0SDSYZ4XaYZk5Ukoq2Dr2b3g
hjIeb1FCWNL34oshrctVga4uZLT7zNyGo7IV075ihiNAWxY5mAPx/j3TBLQJ6+nKMOuTky5S//tZ
V4W1QEthZmiY2wM1wsSTZ9N6pfRsMBa/LlbSMmmBqeMx4VKz8w1q2ePM68q2vX/CMN1ncUV/Eb9h
qLK7dI5rvPaXeYCmHiS07LvArJDPrJrBgYHVXk/Uh6TqABsY7ZW9Za0Ioy5vaxvqjvqctiReWCVS
Y5mUsOmyvBEgCdy96ooBR5NJZYdqpOYtJvYnHU+6a5fOY4sGj22Ke3tXXhLCytYeKn/XDMkhOgDS
BT1Gn+DirNmuYLTSz3FpSSa5lA4CIAJEbIseSlx0xLtrfKC0rG9FXvGLAmaF8Q4c2zaeTErdxOVZ
TG2CxgXsE3ZUHfpVT+cgihx0xGo/MzE0MHmKW7azyTj1kbXxnhJ0qBso4HsXuJF/mWWIlAsgOZr4
iyVF4rorKfen8Eqyst1NQK16VeDT7yfKOkbC91W5Eq/4+pMUBEOuiVv1u0usrtH22Nt3lN7H66l3
IjTJ5rXjWX1+Zq0MO4tMFyB9PUNA558Zrx/85mZKQ2WkYGvvg5eLUJ91xNnwB4jj5vePgLt0Va78
7n0FKhaO2QKzEMxyYcaZnpTP1FyNdufIzy641o6u/bvN6FEuSUTiS+YDPOErpjh00b59rhwob5Vu
mk2K+79IH2PGc8Wx2wPnGUT85sKabEkMThmOGoWYajUZ8n7y0rHQVwWWfaIDmsqq2GLDWHT40uBg
bbupIGl2Ch+Ee5X8sOzEX5M+WeNyxNUHXn99kNSBgYopzUVs7XXrrFtDLD75o5EqaPjuGiwKjSVT
6pCSUReGrB9UNvAAicxwQY0szbXxuw8g7WPxtsKblqxGGJkWSb4seXtwmQMAd6dvqP2vctrkGk2z
FxGRqUUNGG5tsOIYjuJYMSBY+WHi64nti8XlSuLAc0ZvnbHUOje3lCd3Y/HGwAprKSSkXIYKy57V
1xIEVogYXJvH2Huois7PhOdybESh2wWM0pN6NuU5ehCl2g7UauxjUIWGviguZ4ZO9sOqlcR7lFsq
mXkJWdIEfETAGEp+Jd1ChGw3bDJh1sP3nI8jJ+vcNQUshKFAKlpXRfCV2JTJoshp5UleFqKUAAjO
WrUZqiNTR9NF7QJB7LEWm5cOswmcZMw4PpxLFhAzZxKzrVsU6fmK8XHQjCLDTBpzbQn6PNT0V1gY
32tbJTwg35R4fg8XVGO6VXenw0AoN8alhfdqgLM4/AdF/cN50dBgdUZrpKY71Ij3VCAtZcSCxWz2
FGie6UKsH5I6j3iDObtFXG8qLvzrG83KvJVs0eIx5JY/sFxS4L9Qmv1bJLMKVjsNFy5AQwQ/0BYH
2BDAMQAndgsCGurodAcMA5wLRsmac1gi6e5CYo6IXGUjnCiDzSLy8NgmiKxANU7JOiTWpmoTZPRQ
/5JfVpZLLQf39Tqhx0YZp++G++rvR3VuHSZ9Le0S5JLCIGhNZX0IiWX0eUAve3MhZYedsGYC2CeD
goU4xLUMK766v3YFFNZmplmpWpx6lR7kpYiYCEuTUQVcrZuY/m/ljbmSxUvzQma2KSTedexY5UcW
INeOHda7tfCU/TvtmwlMDEjDiljqI+O7NoKN0w9ROIl9w6DrBup8ZUZW+DUEFwA5a8pGMv2ZwuVR
M2p8qhv7R+g3XDtSnJYPSJqHvKWYoYLao9R2+QXCizjCvRCGqWCABc7WyRJrSbQ2vtiB4/7TvwxG
+EqXfyPPPCZSgXtCtGS8QxeJJXfZ6FBw6SU5QyHQ+ZwfdkNHegNNgRKA9rRryzz8beeq+um0dboB
h+4XGGxkf1Dw84qZsAwJGE4yOR5I0Fk86l4d0GmnsdCZqd7+G5FPHScC0UbSQdr6JKFOwQTDWDqN
QcB7zw/EGfCpLuyNveqotkylpfjr2NrMbowzn9OdUyZE8MN4hV4YElT1OPZPW8/mPVhx6dZZ9BRj
KAMdX/28T+YP7iiOTCgUha8LvpdIgJitDEFPWY2QKtFO2/SObVd9inij+mbEfPkqVodrb80m3b6V
WGN9hmlIdI6KA/emp49LJuU0Ffofxi59SqpnAzI3tcFUMia6rTTRRXT/hPmuL6StZOol8tjSDsdQ
kNDZ031efq5I4V6RzKq0Hj+BRJ3qeUMI0BjUFx1fGM61Db8sKUslIeQkyDgALgcc+qE5mCYASnNB
N8MY25KKF9wzgqZ9aIMRXMy2oHXeI06UN/sFvw9AmP6U19bo5GmoEYK9YbaQzQbxN0SssAjNIDAJ
u63B+4Fgx1A4TEPjVs6M5YevhjtrBbTV3ynDHRz018rwYEzR1bR2o8mvZ/vWACEOnBevrQ85QgXq
f0vJq/A1vfuQ13W+azN/0t1jR+kZ2pUvM8tKSTl4S++wIiEEIyf/dZ1vav87qmfYRUDD7QCVBSFS
WohpQ3Y4N8iYu6sbS1GcQ5H8n+Rlv5qZM2ce7ykzwzOjDtoLKXVFmMaQhUv1qyG7kUyRkENUd5W3
itGxo7uyK2IGuxMZOSmfUtmTiRt3AhoHl66d4foe7/Kz3UDWFO9B1HMznqWFXM2dRRCR3lXJslgc
sPDhrIrzhyByiBSK9Kqz7ueLqKZ6LKUNGsbpkqIJT8cyQPbSjOMLJ7kSnHnQD8uYRSI3HwVVOV3D
fTMY2eyeIxf0k6XBWKJpMwpAVtMq2LRO2jJ3sOPcaqvmwZdnJyLIYMaJEWViURhnGqWgco4tuyX2
z8eRAvjl/LBMQzWfynOcNz6/jnvlQxanLXtOvRD8XsS/+lkML5Pf4KqCr2emKVWGv5fYvLpL/w65
5NavFtm4nAItLS6uYBTg/V6dcHFHIoldgUVKH/JpjQkiBzdnRyJdUmg04f8m+0rFWE0eMDN52NHz
0XE4T4vJfRpcqYFm7hRfFjzo2myv2gol6fTMgDxRt8cXqadXqxKfo6kKtSY13y9HFjC9oRteY1qE
ZFVJrRczZldjMwW6VmZovL/tc8nwVlRciK2NMb9elpBc12kxyg5X3aomPrzjE4YK4yq3eArDV4gz
8OP+z0w0NhGcQUCZmoaH1jukRv9c0lJbY+YbX6xbE5wkGwYHUBCaWSSZ+76ZcyyBUXw7l7mU2X3l
nEMa+LtaMk85ZmCcvHcz1Nm/KRbQCIx9uT2d0fA8PMkLak3ims5RRaGU4Z/siHfeX2UYw5/w9+WE
fO0cA1ufo7BwcjRKQHYju3eRLiFyg/p8fF1iW9zxj6++rYxVfIIkE/8At9SoYLfJqxpmJ/A6G5HD
Tib84uavfOQ5GX+Fm1rQYBaqtPV4nVmf6TJKw3Phx0KFzAE9pfZCZqxr83VQyP9plH6uQ51oUXIS
cAfjL8kp2AQ/TXjuK7EGC8fznKWWjzJFojxOA3GO0bv5pGsAaTiJe0xq8UCW6dTlqowKjMAWbhMF
zcvWuGC8dXyCOO1vRONnQSJ/JUbyi+0TBPs4CrUdn1vTgMh1LqLIKH3f+03MifodgvlzeYsut76g
77PqZLqZryCRQsmhOPlO0IkpSGbhvLryRq31aA8+rKub4CwRVteDgnuzGu6VSEy5Hjbb685iw0Uf
EVB2oAXXvwqkv9yGypN9GEiBGPZ66zRpPQJe8j5Q+xJSYQ8cQK06MUG4hmGZxlw4/kwmUPCRUuRJ
axxQncrSfGqwzxZcU8HQJq+CnOhiOGILPL57+jiXZSv9y4+WcvMvDGaEzQzgyKTsqF829/+AJOL2
UmEdFxzde6Foa5mEXhiks4QufWzOIa8x1IM8wmQJTBOaMbVob0CESbhRiK1w7qq9dtesMv+yBxd/
fJDLM8bMA7QZUeI+y1jDMbcA+XP3VTvi8aZjU8FTU4DOV8Gmyx0RjFqqwLdg0wGWttrPACaaqXy+
4RdanLRmFIG3gsKbeK8bdO66x5JbnK6j7yIuApMzLUMhgwT+Vq1KMZ7MkMRJPUecM1P0IRQPn9wF
M/cbvg9svm1F93Q7SFlAnNu/sbGecdPPg8n8+MUxv0VKJDXLfujxOox3R3C9J8QDGZHXpky6GrcF
Me7/wWPt6lHELw/K3ax1NzPRHFE/uSttAlQ+U91uZOjM9qhMGGv+jpZaM9GQNWkG9vyQabvOQmFf
AagUFJ2g4XfWByAxcxRU49wxnFZZEYl9TYo5prsOiNImribLvJVuhn/KIg0DRLzPsziCg+hkiT8T
FNvJYjZKMCqgtlr8wV/uHhkGt8KN7KEdb9VVU5QNcX3tup15mx00FUpHm3EOKvbNpPUVn36aj16+
CJcRFKf2koW4m3dxzkhXVt4OLvI7KjUBpa0GIerfIQylWTCrrLrGWssxZnTeNrCUINl6fWDZp1xu
I1rPMgt/mtxGGJZldkUnuSNrcA4UzzAAcVS1nRpwh8gceXEMGBHi1Kw7791peOwJ07lyiaPlX8J2
vdH27a3TCF9sX6Qs+jkDEmYphqhUWEWdMlkhHGJrREJ11+qRMHWVpHb05pprdqvl4EwvCl5PfAj3
5IEFcwlGfitm9CSqPwkQyvPhkMFOoG6LQujdXgB24nqnZ/2/M6ign+h4xpr9E1xILa/7MBZsmyh9
AJzn2hmATOwBTRvrxFsFiBAoei9qvi+Y0++uZ1ET/kdXfOgclBbimVG6n11IW1iRNvfpRyF9/Pim
FZtIO3tvGSGEhnxl1s64TooGtzb/NkOn8Efav4/OJzK/TSzk9rQOJwx6Tjwv02TMv9p2zAQkWl29
pBvc/AtiZWHoGXgdSSD3SFVr0ieqbjjUVxZE2zFvjAbWYNl9nWqv5EnIfyXQCZzU95LNKmKokqqQ
AtPP+n7PwWklfbAjBzut2St8TKm/RLTSEGzyaYDR0WMi4k4sajxOnQWPhA3l7qK8vfroqp2ZMvFY
XZv/8gztHAdGQCMZQSLsGjmk1XOtTiehT7hNCFd7nSVqPPJmUwH75eFrv90jdPUlqAQolYMIvPev
1H5lePDqYYwgR8wc5W8PVjByjB/3L+OcPyhb5tYkgoA5KR8g4yGyW5Bme7zWWri+HBnAzDiUM2Vw
a+xd85wwVyOGnUqCUdEkc33vpcuKZc2xMNm4U6B5M2YTPH8Zhw6R77f3LobDZjsEZ7kuY8xrDpn6
FqlHFr04Hs2jlkOySrSsdj18LvEKkqJUa9qSD2pfbPJKR7luLTwLPQoNwgHlkosat7F8GqmzTUSs
z5Sf8xqSuJMtJYxMgvKeAtH5slppHBwJSPXFRXXp9W44RGa3a0yvIg3seN59Yi45K1AaEpJw3ixA
X+kp/ojLjSQucC+Uga1Ooq3pXxOEYo8+wCa+hfjJV2j3cCiDYBDBcaTwL5MtIOMogRQfPlq7B2fF
KRbC4EqDGfrlXWmVwuImB+MeWL6aGk92VNwPZ94WbHCvm9vqKQuHJwBLzG1G55WohA1UeSGMEqQ+
k6pdRVsS3wYew5TcxpV3cKnP8S4xewCPNM5Sa6nIZ704bMuMzVDSYslFXEK1YiokQjyIGkmF9Noy
X0wQoirdk3oAN9/ap/ZU1RcjeE+eEs+34nl3fGESaNsrzHVUOvJFKo4Aoh17I+VNawEQGOEL0HAQ
b23nf3ZLiVrorBIp5MqayHoaLzYDLeQJjNKm9YX9BCqlG+uMZ3C5xgFx8PNioC6fVLpcSllSrCYn
PbJs781tbuAjNp+STrd8BmqzoFlSrArPZhxfDpdQxxtL0JlV8u7fA81kSp95Gi2B/TH8cN3sAa/T
VC2rPlc9PvbYXhVb2HL2XXWIILhZvnvOSln+FZREO7b7X4T9sjLea6Er8hz+bajL5PHiG5ubNETj
ZYShd8u+uvtj7fLs34/99Od2lcpXl3TXls7tYqqK7IBVfClBRLp7vT0HSUu7MQaf3bwho+pFrtpD
bCBcgW0KM4ibBNIkxclFo0K5MC8QswUJ9V9ygVSpvkhQyb59hQkiwJfKi5Pe8VpNnizvTMM7bLKN
CPALtKZfMgP0sMDePhz50lTUcdelvzpHjDj+qXn2l9cpZCJwZuWmGKA566ulhZu21bKcQOiUVXH7
+JvIfPAN2SX9JcWO2pz6O7xe3y1eTkmEniyZJ6dvWye331oAIKYPwd196N8MM1x/LDd4FUAAxPuf
duuxcE35pdezSZTEuVhOKEWP1d6MPFr7EKI2DHGhh0X7yVmjgHfk9NvU4+CL39FWG0bjUePB2h1Q
lQHEmjxN7+P/KaoulAzcTXAMwCUTHh8IMyHkF0oY+jwvFaotP5kqP3dsXAx6V5Hz3JoKyKjsU0HU
5DxGD3SSVUuo8bm9/TEZ69yQVEfZsckGkIzhxrhYKVOAMVQaTo9+uankEsyowAy05OasNi2wi3Yq
9Xzxz+XGW+AB/1wZLrrOsQyyYWK6c+PS5wJs7Mcejyt3cD0HvIw+KGvYeaEfjBywMwjMqwCaO6L8
miDXf0Zfk/q+sDSJQ3lo0JCZDUHYV2gsktrSv0VADG0N7KGleIvW13/43StCEIYzKkWj6BB6AgeO
ZTEXjzmeIhKUnR+rr6PV3oCpl2ubWHhjcZT4pGWI6yO4qIbT12vfufpSiPj3uN0dUpawUGgdeffU
+VHnxY/3Xaepl7HeVn5gMEVAsUGjUMZhYHrZqfnnKJV8A/3ZCora6U59AamwPVTx12DWn5ZGgnqc
gBxppXnCC2UxJaoUG2Db1o7AthKnGxudsu8WaoL2SiQeM1YVgl1uGM56FDWCD2XPa7kpqDGU+dE5
weinGG8EoSyeuvBmMr1t/6n2SfAwMoB9V/2di0+R+ZuZ2sXg6wjBAWZA5koa8EUDE1NKwdceSfCq
Y1Z5DEm1HGsbK1a0g13BFPfBXmsdilWHYX1R4H5AEwNTTiXXknWuwhM8U8qE4QNpRNsO3e6pVCnz
TUKZsYvHms64UVeffThczXkuGMjk6Lllq1ImY4zeQdw1DdkLJ8PlZeLQPc0IAwdVcK4CP3VIW/4y
TlksZibBy1pYe9jug6dTgX5ExxZKKZC7zsSixTisAOx4CKmDgyGk10pRBQQTGyGQJMDrzBaPif9m
7CGOxLZF2tizmzlsvNcErgMbzDzi0F7H/uO63o+DEOfzf5bIWuN011AZD7hzrddNvoDUMtuP7kvX
vjb06b/aztXHg2veb5Fegsldjo5FXXipic3iiqancAwJIROywCIUgmXxdAqOOP6ZFU0+EdAvC1iV
arrGJmuhESHII+JAje6oTTQWZWpRhqDJDicbAZZnDlCGQm4Tz19CwRiHLGzi9/NRmh8TtdUnemnQ
D7G8GEFuKnh8SHlSekR6p7ekoIhpVFLjA9+pJruwqS9F3o0B6mIP0i0h+AxpbsF7azm9RPs3L5YL
rCnEie11XKDNxn1b0pDmiM179XmZwFWmSQdMMqYKZI0/CnXSqJsulklPi5vqzblCleUzj/aJ8yfC
1rQ6BGcs+PHvEAolp2ZvzPq/dSERvDKq/AVql1p5bO6pKZyrt+CEn7kwXMUPMPWRD1qm8DbvcxBE
WqJKxDThCoj5N7NNaxJ9zEakyz0VWwi/dlk9Trb6jRiBP3HvOlOHXbXDlpLSh3/MB3yDtpB7/6J5
wp4dE31xSXUyWVcujEG8IHh5/O7MhOIMsCWvrcTkl2FWfwqUkUix3drn2AI9oaYUJLC6uZVl2Qrz
hEt3VuFCgDoY2bXXFfeqPk3BiPAseArH9W2HOvMjZY/j176Tb+S+XFNS82yIVWMo1pN6cK0dEDHh
0VriDXKmWYcwS3al/1FG7WJYesw0RZM/WlsEwRy1V4AAGFLbZvFzZL9P1OhzIvK+KXYbgP6Hkeek
TqMI5YEl8HG91eaxG4Awvv+cejD1nXEQNPIK6jElw3/Gz8JR+4CwfBMsL3IzsTHc0Gk2XKD3MA4O
eDjVWcEXystLQfVd/RyEVskxZn3u3A678BMjzy6Io2DgftscudP5oGviUURnWcV5BIV2qIkoC5V7
TifTWl5Z+WJ2xwWc2W3XPTudHDsvRXM4yW2C9RqXxMkxQ7JEaWvH6+Wl0YzQu1Gs6fzyL4oKnFIL
AIstfXJCy/tRhRS3Vt1R+3Enkw+RkuqbR5tQAqv2Dt+Qdp9kbpAr3NI7e3MBj5oB/4yFBTMncsvt
/+a51ukgFZ4kTgJ4alHcvfkVQpyU9gHJehGN+fMN/3600Hkssz+tFE11psC8zB4X/aghGi5No1F2
FtAez1KrnpOFD4rHKQWr1j3LEMdUHbmqtd+7Qj/9V8lS99JpsTGse1nxX3a4w+S76ojXObxraKWe
QvKwrmXfrhF1hObkPqrZypqw2ug9lHO/1tmF7U4Jf4iTaaOBCAoXlMMb86bUfjhHNfI6v46wLASl
BhsZs4MaiZKYez64gIgS72yMWqLGwGstXtDGA5uL/IyXnM4uELkkuxMCq01OPTWlLuAd+r7TY+zy
yt601jnadvErYkH7pTqTBf/qKZkeNQJoRPMBC4fKGxgZ7AzOVb5OtZNkHvWmB+4DX9eHf8IghEn5
0fg+WIl9Ik0sLDkYxAx3DwO4I2yRGZNKCgZ2tuhacaQ10Xnh7dhND6GunTjtzVtNuQWW75dRyy4+
7vFDKbBCChLyB2OR9VTbnhfS3ITlp4ahIG5htzjia7gAtI9t0FuKxXkn6gioSOGYx15YM034DuD9
3BIVROpqzkh5muWnHoi9x5pDTO52R8XdGZRWNDwhBg361KfnN77iL5cneyUBcrq3uUh5SsKm8yk+
xuzgXzlBINNGXxxL/T+2j9Arhe2FsVEVmrnbtmLWSCj5+OhQ0Pj1GDut0T2NFYri0XF0Ns7ogCTB
30hZBf1ZNiZfDj4jSTy+CiWFP1keFCxwD01H8UqATAVWjX3YDeXg1Thmat8D9o5ulUYrpYdhZNAi
NFiOlPqomDgKaEQlBA0njyTRbi5QxrwtJV+2NwFnsGLf3qM0SWffHQbdCeZ3KIeReKffN3/e3bRK
wytpgpzOVl8gFVUib80Yf9Yh0SfpddY3Xp8QtaXpHQlDlk9sZVcmSFI9pcK6F3i5oneD8d68h9xs
xJUn4vkKDw31IKWfVSm2XKRGamLyLoHpGqIIcS42u8298LzwAmq8ZIY/rQL3Ue2ZimkqwIQ3D8i5
DL+R4O5PpKuKX/ojNCE3Z0L6soj5DQk0670FTQbRCn5tAv631Bv/3FBN26lbg2guDp0rw/1hTgrn
sOoBPQuQcYCQNKr1VMLg5Fd7Bbrf7rJA67++H4RSMhrFPV3XM3eAKBifTfjXIwcogrq+64PUdbyL
xnvnYe2TGiHYGunM7g8WZTXeltikzMJ5O1G7DpS0Jm2oiMq4kU7tpzRJRJm4D8Vy/YfMhdl7UKes
B7FxLD4eETbeURtKZLVt6X7M5U0rTZj2hYk6MAUjPJhbNmGycqgMS+Ur6Ie/TU9CqlJrmqtQLHnz
yuMXCG6jCECs/fxxow6enn5dgmP9YCLU3fSGPdqfQ/mgsz5nK7cIqAtBXg1gnIlOR8opgt+48eP+
risQR5VmQVGUtdethL2xInhfbS99rqpKVjOOwCM6mIA4jNvtQbv46XERjbbRmZMv+ts01zFelNyS
++3ICmTpPIvUhaFJQI+7gsNC9MLhUcVr5cKsoBwWd9rkbeny8MpwXA1xhEL0wV4e54MyylOx8bzX
xGx9TLNLGc1wp7mPQf3ZmG7OUCuP/9l6Vnb7LGIxt3ueTX843bSlTSJfYaEBwQFbJhgB0/ak2SOT
CwtQnVRBGsa26FkmncgM9bpeeNSAJknCxCnoJnrenU8TGJgx5/GKN2WCRiPKcjdTRQiIKMMUVOzP
C17FHSGLGIooUITdDPNUg7o4PS4rDgh8mYfHuNEdFdLdqE072t4xA/PLaNFGrY4Abu0ojcczTxFF
B2o8uXUnY5JLzziO0L4wZHo2vshwxBXHWDLjAW2HTxz4zW04C5QEiD3INYT2KpyYibJ7lgy+bAS6
bGOAESU3S4+cUZO+yfGKb2dLsABwDFglAiCSifYNYdlnpFPME9ZX5JaHeIl9Gpf67dXi46B+4ww+
kV2uqAhc0BcFujAR//niU+daaYZ8E/PnL4vExDH3ntwrPCv3WwVJihASxAMMpz+CKl/cEmAQKbAv
m9CW5+Bj7LbBqnKjClWoe87CzJ0vylCngnoRdQ5HAvZHAvvTkhKR256J7B8WGmI0IfuZolCnfp1k
hp8EiaHQepZo4wodSFLEVOxoof5Yx7H8Pdt18E+rauelx8YvwvhFXg9t1kqhMAlxpV4RDi32RMIY
Dy1safIwm2GK84DNH8tiVUHzFEPm61mde/IFvF8rE3ZSKI5rHmTP2m3681SBcOTKtCB+Zb8KF3vG
aWiOM5cpVmS0ZiHEF+XIcziubib0twP2U17CJSyLytmFcAisT3mmx8YIhhrKCnVNlSL3T6Stbmjm
lIkAQUaRJUaM4JFKKvZJUcVade/Eo5BJNiX7eSgIAUGi8U5mqripIy5nvl7gNykZ+9HSs627AO8o
uFexgdVbo3dhWbzDED78dyPAJkx6Kq0XROflAJJtib2tCwvD34czRZwfOdKXXkWxk3umlHy3+Ktb
TS7+Fhs4wSSFSE8C599cBwSF7R8P/V4sT41EKTCf4l/fysda8NNJpbV6YKXoeAi2PHg4bhgW7+aO
BI2KKdhhVCzePd/8zPo5CkqEVB+MPl3CZPmbyBj5LBApvT51lunE6muZxcJYV9Ei7K3GOzKG0kr0
FNu4kaj+f01xqH4Y70OiExwNA9kdGa8uBEVHPabAijlHL+VCezm35dpmMDLs7R98ZESDowAZ8rst
kWDptgh/7G9RYMMo/XL11FLOZ4KuwnRnd0ifWrSldZCs+rGuZp1dJmYPj+mCBYoI4It/8QjE2Gzy
hxQa97ctwcDCUklCgAwzZelqLr8VEozciH0QUJS0tuqlBi8heTaRcMVhfgIRweqOuAHKp8EFmjZH
Xdt1IovFsCOPE18pp7A0djx0Nu+sjdDUr67sI+f27GYjQc6VZQIXJKzyyCFpylQpGJcYco4bSA8H
+0NpiRs/4YyT5tEFZaJeKd6ORwynaGhQZZWn3990n1kHguKLmY7OXVGQV/l7vWIIsjPY6V6HwZ3W
hniYYhjA/bxvRuUo53t6+vwe4uEb/kxaTj7bix5jI7gzwKHPZsWDVkB2MOyAYVLT9D6fgVAKyUWS
HPz1Zt2KevkSIb0KBNSsYRSfh37yGbiOwoxMmASzcNekjvNkdoa28fBpBFjl9P2g1YYE8oOxzxDR
U6z0fueM+Ik8FlLAVfsfUX46l2Hz8OZLXAePszofGMt/1xR47LOVxblTAnNxdJnkMMvTVDBUVhcD
9eIGTXl/l0IXFoRIX0G2e3cIKJeR+Y77fi3KMQbJAA2UOvRs0VYKmhYoJLoTm6JcuUergk6vEOYc
tS0zrXUu9y/40vNpgYrq+q51SFjyVvJdPEPjDvaMA/UBARJjirgDkOwkbs9eG85BcrgVT7UeaPOa
QFEAH/UqVFDKJj8sYj1hQpMOs5Y8JfKRzex4qqBdUiXWkAeqtwIMP/IMlx5DO7i050oysxcg5JRi
ikjDHSRoH6k2kgaRgE7DpHkhFuzphABxJGe/HKmNB/5qdchY03iHglJOZhe7OS36UnLnnnz/NzuY
ocUtQUBD2Q0u6fGOjZTmpfbFVftbFBXASuiJGklXPtapA8BJk6QchdTC5KuzY6rro5Jb3ozY0yGz
59Hcyq6RlcfvYcmpu52SETDRVPJxbhNi3y52FTEAPzczs/vQN9xavjJJSDHkQJmKaJGShh0R/zGu
HhuEDD6BZc7wvmeRJMFXhn+NpEszabxEDm9IOljor947gAox94IC7Wwp8Rvx6XBhKQ+JeSXtsTEV
yOQ6p3WTy+qiXMESU07+nKHl2/tRDmDARMexzq9mmyoLDSc6IoJ5sj6JhzkuNBewpFcklrUdhO7d
r0IR+w7MNQ2hETHgckw9ZPQ7R4JPXswx+EWidtTiyF42NeIvUBK9MuJGtORegkztqSNrCXzdNk/n
+kwntYpaQpuaQ/Ucsm9IBEGBfSgZ9zcpRL35qynVqD+uEinwk6oWSPLIZmDHZhhn5wdhKwCcT1X6
4DKInqwNonmkcqVpBqyPNqgs2GJNTLCWIUDC+wJTISMV/Fum30VTVRdPDtTwM7PV97w3pU4nBYIw
qHSKCF6FJ+nf7K3nJayCn51KqndSgxA+hSY1BIKN3FWy7L9IShwLfxMsfYEngWwsc7qhzy9vVuvl
Py0F6sWEtndU6SxzuG4cxJk8jXZDkKyKM906QOV7jOZL71+6gPOBQ5CP6SwFedCUdbweSV2SGbJS
boDkZUzTb8U0H6naI3AocM5nifnMBDJgNMXkCpFdg9aF14plQs10YcwdK9sIIT0T3SmY5M4Wwy1I
Yp4j1CgPtQGLe3unZDumYVqfgR48lEO+/WY9MjKnRgfd7tOABN6RRQnEzqSXRxOe0Q44x6N+gpSa
V/w6/GJfYB/QmCaJZEHCa2+p8edq4Umr1W763cQii+ZDSRbLpaD1z8M20huhdf+U5OgYV/6U87IY
p1emwNAuDkj22U5RAFlV/TE0pRM7WGie8U8bKHSVnAGNg6c+dCFtsuQ+C7NwruAuXhI+CORicB8I
qPo+/8p3+7t9tp0whhP2ssx77DnAzwpx3+xFWEkSv6cZThZWz+FqgxK5LozaLRhb1SEfRQvGdOxP
lU6QxK1lbS6/T4/ZbUKqs8qP2vV8GKQglGJsgsbCokd4Jh+Zu4WXhUttxIFNpO2hNilDa505GxSN
lH25BRq1bqXHHHmzeXnWbNyo1xHPFySzgaPtNKL1F6fOnkJEwlZ3kLldZJ8FjpMHL9DxhDIjE5fG
MjfGZ5PMwvzhu6Ln5QAN+ECVg6xDoXw2rtioyay3+fNG4wQVd3MMf6TNsQvqs551PIOMAFxPiakA
/TWT3QhRHviZW57rot4Mwxp7olrcCuPlgx9N8QeSIdzR2ZrZ0wcTaWcmupTVOQzkyfBeYeuoMmIp
22y9by6QgAV2vXnFRzqBZ2mvklUnwbrQ27Hnh9XF2GintYhheidwpw0bgbPKJLbEuv8mUjAOoEAX
dEEuDDzyyOzZyEeSUOeHy+v3bsyJwDg8mGUgHjjRZVO0xMF8p8ZmEY3unzAahgVgUwA7NpKgF2aT
H1J9Vryl2OFxxVPUuccw48g92uRxvmEJg2FXT/va7wQ5A03nZSYmR2D+yvySyXfe9tDoXeECIqvw
JM9i0cyiemjDua8Hk6tzaiSt1ipbqe0MjnV+R3McwO111BvkxsrGnWwKu5wbiYg7grQ1/pGp/9W0
G+Rb0M8R8PjU7QmfkGjGub5zj/ticDE0n8Tpzmt1jQtJV2Y7IB2gW+LPE93KpoNk3525LPZeGPhz
a3VJhl0B6WRTX4DXNy42yew+aVLP1S9YI8/fOKptmGos219tUtLxNeez4vF5l97eXbFaw8PJvYWT
a3Zw/F8igbbgpEvdVFFea06SgjQ+BA/945eDorlny31hpN29tXc1liMTfFh1KSRcF3+Dhujv/QBb
GKMw2FU6n38qvlVqLAtj3wxYlrDndQZ4nzebQgSiJu/DvLZv+UC6I9nsYBxHAA/cKC6/KHtRy62M
vgSAOoEuUiFT1a1SXNSbyfEw2i33mrVi8gArTdMxTxtguUP3EJVKhjPCsEqY3r8rFncj0x9BKpQk
smg8TBYs8QlSEQ+f3sNV2Ug25UDvP3VGSDqJUBeLVjEm6FxOp+SvJm8bB3oSxo83sZySoU+TBc3h
ooYreiKdQHxI9XKxZcuHx8zgXJNovKtR6vOEhqqaFTruAHfX9BsG4AzVE6kB0BBkYTzbmm/qvLh5
qa8L3Sl49f/Fp+iPXj+oRtB98cJka99xVQ+Mcbf0cOT0oI8yoemjAFTBaEffjzi6JOu9h9N6VR9U
Xw9bdm/Bz94DBtcdCwayNMi2RkKVwYBM69AIPDr30FRcQcXmR4SCQ7SojuPls/uuQm8ARJbw/lsf
tyzGdqMuaXav56+54Cx43tJTb3NnWCw+7J16dHqXaeWSQBIkaMdJstEjzQySwV9JNFxjwk/gmfN/
hIN1n20oOeoeOGTV2tnhJZ2R3bTDr5bNXvpgwV2luRCdg4FE1qgj3hj4WZ6AvVPgMPr1skLxhrSW
pL7z7CuS8Jgg3of/RmOQaOtVz47ytAiIf/bLiwUGkxwPT+0ezc5oY0Riqgv7iYQnOi3NRpbvZxJg
pDkHYiXlSEMOW9Gg01/6I5wNAiuCif7X6pgd4WDXyb3831HG7c92jKQ6zsid/4AZWBDyoV32ntf0
F+fiZKEkfpAi7PUAJnQb8Y/GdwgsJx/EJdwy5+y9vaJbJY8jl89G6a5p8QGFFwvjEoZxxi0FsnLB
O7GWRApBuuWK2KUUn7DpmevwTOXyVcgl5rXZAgnx8UlL8X2cBQAl3iOll10hcZnSuvc9mLi1Vxax
1ZGq7ld9dxeRh+psLnI751su/Y93uvx6nJZUMQSq5X0ckVVeYHxRJPRxdb8SF49f+YPdXWWwsWiZ
ZgXd39qH5eyRPIX1AlCWwb+h+veFhir7nUVc5tShU7TVwKdfGEfxh29Rpvnbxw89GTQxvgsjVbdL
FEt/c+ZRjBUt+q6+npMamqK4PFO+BztwOFEmjoQwY7kx/VDb1aFSMAqsJKPISdiNhFK4kNUheYHU
7PcYzv2bSEiA+F46iaLl0f2f99+U+7rTn0mpW/yTYLyWTXb4EQsH71n2TuHLYvm6UttkIuy1FL7r
TnnSDmH1hfd32+LetrIfKGEXt8UJtbILAQK81VZASrqdpWtUWlVoSN5z15gVXNYKcXQrPRcLYeMS
z7c1yoxDYD8NVAtskHS3ExcxhC4B7NjAUvshvvDSuFiNuXvwKa0CunsTwLFn5kYVtuT1b1GIvfHK
QMQT4GYIDktXyEbpRtRcWCoQKhe/HcPmNaF6pB7UUuyKy/YtEZgVYq8cBLwHdVILkPBqzRoURcoe
zgJX2BfL7vkwFHzdsWgJQb/R54fexqP3/KjBFjDJuwoCc7EZ1hn0LrBliwQhIblLJEcUCOg5OIou
AS4mf+QK4Y/cDSwR9zbmuVy6m6zRY3okxjiKkVAoxhryRVI3aEFe+0dl1iW7gxyXtEerLgwPrXSZ
lDvuWjnbNxc2Wq/cmFK0B3FrBhc9ImJ38P+soV+CKsR7OKnxRxC17ZHUry3uwBEQx0oYpLVS/QMo
BBj7xrpN/rz/qz9vtsBc7W11zAZe5XPDd7GR+hBPOV2KqLo0dN5cYyOkGYEE5fmuO5phWLY9BKHZ
fXPtHbG5MbEkZ44bRctRSl2cP3PCGHZfk+1ejNTfeW8+VlmjKNaKIubGfb7AbVaTWvaK1UolsI2/
yOomDatxYxTuaRtdwhNiG6ziyZc5EIBU1jMp4g05FdRqCLfX7POjdp2TNsuxTXXzOsIg4OsTp/GL
rY/s1zUY0/yYEhRHBk0BqH7WxfAdFMCR0hfiPf6tr1q5a6BwK+hLMEYk/uX+xB1TjQMXJsnef/sl
H72tYX3/BN+oYKATAUW5ZDQmhCRv0dpmt91moYyQ2YGWUrouyz+6HBHCoF+0tPrkQZOA8Wb11JXr
+6+Kfu4nzb2u80H630Q7r9q5lfPKU0WzGnLuFAgK2wFTdjt+zLSZQUFafoLJeuLbliB3MjZ/NzBU
qI7u0UhIlkdJhCj9N/2iqGZ2gtY0OkrQHCp23sWQByKdgP7nCdhRzj/tSLDyx3+/xU+gl/wsioxH
h47c4F2gjyDsgLTdXlFQRYVrSZXrN7lekA4Fa5yNUPbeeCTPS/xOEyjv4zkex8FjDpxyK7UQIaWw
3+SEyGGgkQJm7bCJuW4C+FKk5AH30hEAStly6hHAzfFrPg+KX4jdouMFkaTvYwITqfL/ZcJrthJB
OciZVZmNxD+aNz8QgHq7+3sejTlgqH7azMiQdEPv5bBqEPX+X0oy5AaeUUBvQvgx5HWK7+cvNPcz
35XkxVmfOQttXL8O2sR9lGFP0R01zSDNLjGJylRRFhUpRefC0oegpRqoggH/zGZ0ciFB7J5HeZHv
JLxbt82OPiIaza7JCTE/1G/UQ119GDStytaHUxoMZF8TLa0WV8GMruKFBwnpLCAHVEXtQZHklJlg
Zjl1oMVbUWxSZqgGhD7WX1wxcP2VT0wEACSCc4IgbxBGkDG/0ts92eeA4AhzGXYYXJIDxdhDPrh3
mzs7h+h5qxJKMK8GTWNewLqnCIBY37m1HsQ02RwuA1LkjOCJeKvDdkw9XkcH7NVa89MStYZ/1DLg
9KjTbfy8Mk+JI2BMOnrspL1Nk39su1bho2TzLo2td4VI9rrCgD3dhb7L75eyPenJ/6BZ9Af5zsi5
lOUGyn3Mi+Vb6bpwAbrrjefG77leq/t6h7bgOeJp+FAIb/h+rN5GBJFquX6bgZN9/2WtbxLiOjcY
0H+/0jbnaq48hmH6AAekYE92iW6tCThKrSD/mnuaWXA5oV8sF/C31W7WuqZCGYxGMsvT/u/h55pW
DNh/RG2qIHO/Kzw+f6N3cJj/5pOH7zzRV22HRFHReoIqfbuokWD4Uh1pUYempoAtOpgd3FH7I7aU
1iao1FVO4xTJEckBmoE+yVQHFHtTbLK2FBJXx/OWDZ3Vj++oDu15jhV40ZUa5B0idDelhlZXiBuu
G3Yj+vLffMpyJzE9HO9k8KYPouHi4V6ueAK+4gYFEeeRhETSkHxWTYeS9tBPofohmXoZNcIHt80Z
gS9iyxJ+Sf9z6dy2dSrZpoojl60K+tV0r5nL32tBjsbkv8EjfJAiaUKlNjnOQXLXhExOtkxvplDS
5slD0Q3CvcmwXbAu6A2bxGd6tr6O/oLfTqStRrYm7wP+UsGYSxAMdeyx5sy+gfVnrgBiBW5Gotcg
uk22UdQo3wdWOXFAKFgCPLrVSOWSAmHnAWYPmj5GEjtjHRaZiaA6ns/1u20VMFCyfCFW3Ci3vr4X
ZBYhHRSRbr/HA+n4a+HQ1SJ9oEuY/2emZytjtRkNHXqycxC3Ci8PFAUJZLKReUjnj9kvph9zkYtt
VLemje0I7Ncmm2g4Oc2GvEu3oZuePRpteK1vPmNPra2K4Pir8DU7hCf8QhWboejjpz09wdgB2Tps
jSbm+qjR0qiE1gPgRyfbAz8fLPkwO6l6YtyUIM7mG0lLzlCdmfsb2aWO8leYerZK2JE5rHDOs958
OjDHNlBTVgVYnEX0q/7D0KbbuDB1yATCp1yQSK1vSIQY/uftXQXDvaQh/uf7kXRM/cMg5D+WEHqR
CzktyVz3IzOKSezGVf8B6594lcEY655m6FCkKfL7Sz52GPzGzSiWhZEbmYEPcvI8GqprAPn2J8NZ
kiWxoPG/g/YCxO+ilZXj0yCUGSF1IjIN6bhnB45SI0c4lnvoSGzRsWaQEt7ln8lTei1UBxT5Og06
pP+DBoPehKjbHMBTK9fOyr3BXyspWc7fty8CtrynsGBz/Be6qw8fV2Fr5ckJPV7tadAJFh31l6Aj
MKlJfO5sugSl542HQAAoE48htRWMetQJzhvwCzl5hTXVstUyOaAc+SZfiV52WGrsJ8Ilc8FpIIbH
YbGIljbiDN5FcJnN9e/uvy03CeowH8EMK2B/Y3CW9IYQ7EnhgAyn2WYXjq+fH45d2IK8mbIrpTC3
hvaq1cIvcpOCGBs/mgAsAd4x8r3o/vH6OzDBRvTbFnsiQyn02Xvn248gfW2a4grV+EMhIJ0/vRks
9aXlTCNMn2iVIjybE1ccA476TtJBk6pPuXajF7f5hQcaMCNZ5N3JoHP0/HgLIpAePSSz5RrrTzVY
4hODzXd0pDEzOW1CDuis62tufrP+Ql4Ip7m+rmBVm7IZxYE+u7P4LIA2Wc3sbK4EsJV3p5m4FBSJ
ZZw2J+BbwI1n6MFEQhKgR6k4VV+voqukDXww/hC3HqIGn+gPx8agPEujLmaWxS3kj74ZcSGBv5VG
jG+JJi2Y0oClxGIm5FFBAsaON5hJz4XKUfXPUrGRoGQxOGoYf+3y9TdGJu1OhDDm1j4aCz99sAa5
D89VDjHO2hqXWbZwyxpt59wVw8Jtib7txxFDbWiEQBrsI4x/aWhh+j7CxiZhTzoYxGrVlGHwRl2p
xfg1ynhLv/H9tgN5eA3DXzEvmWn44D/dMLH5wIFz2E3JyGCC8eAQHWHCEQHYAGHEZLHhcnZ4XIPg
NsBf+M7OzQAfI1AuXYTMJyZRnhsamGyH7Vj1+mcVIb1pzD35pS7wdEYtEHpc3JUxFVJLdOkNRQ1p
MM/Iw93NBzBe3mCQWsendgjrtDfhJhx97xFrMEhMtHBariMWr+1qSVaJ/kD8aIgJhV/yl6zTR8fK
H6uukzV0ZisjHYwDO7YxsbTxWOw378vh37i0l0ESSMrTSAxPFc0MD1LavjI1LV7d7Ay3pNM2y6o3
C90aOeBbMH00mN43OAhVH8rzLG3lEDxfAU9McSQq51mHpNlchORguZ+CaMhDZ8k0/4qWEtwWI44h
4PkDCeyTxIvsdMNRum+Cjy1WhUnFilB2an7CDREJsapepmYgi1lpRbIRVVTlCz0erXRvhANV0FTq
Th1a5Feh7IeGiLVBbsTBLSXuSGCafRBmlnCOt7QcUEfY7lROwMXWA8P9JChPp6pucUoXx9Ewhywa
Hwb8Yabs3wW8gVPYi9pnQQhUjDnBDuLzIPldWjXPvpw+dblh/IpBtIc2Emlm0E6rhpE58v+WXCIu
r4gGHsos48WcO1OZZxfslyGdn6pybi2TW8AdRq6e+TcNAaLWdsAmk17eiOOqDBH3Wkt9RoUrVY5q
PuW/TvPVGMGsjh7XoDxNPXiwIwHnEG6yOJAaj/1v6QEgemMkxx0/ZeDEdJAT3eMUGbIHJPzGjn7m
JgM8nTvMQlxRnkSZgZpw1IaNS2jTPIlN73aNq2HTZjErYijX8fenApDJn/IxDajXKmInejC1DzM2
57uNYW8K0u9btJR42fyPmx3dWdCHJrKmy6kz90b0pAeEIxc7eKO8nS34dl558CHGZmKM9aIDbZDe
BEoPxI/Uo5GMPhPZQyk63TvGNGfvVhUj0d01rXa02Z7rlF6FzPvlsZSTdvDpTB9cHArzlemmN0Co
BnGa+YfN/tu89SI5bsHUuDGFZVzwDfL+W5GSuqHnR3RaRbTcEWLqUOLb/57GDigGvrGtIhWRIpw4
b0bysYt6JShgzFHwPpz1P1/k/iPGto2AreiPzpCEZs7huylPrSO5tnPn1BMOaqPpbs2peaHpq6E2
GOAnQCxP9ZrOTPcTkmr2fOzptC3Cdew76MEgeiMmIoaEWn4kPl4TMrr6m0nuQFXhEuzvTM8z+hbj
ED5cJj7rbDtZlMO4ztixnES8O+vvNCiPlH2WaHFTBIOZF2K8EZFxW2wMKsp88oCvsQYK2hIl1/CT
QQEKhLUbjjW+DfaQ+zDdBLohl6K4Z3SuxCxijVCKDbkPOxL15TmnKquZ+q0cVAj/RVpko/kgLVCM
j1yRq4JzeLb0SB+Vu69Ds9HjOP5WgTHoUzsekhSlWlSkOA44J3/iCvI0XlOw0iBxsbfcc0cEv59/
kOHWMWZp0+wd5mlCbhpEo694kQR5grsImGX8xXjew7is8v9+fx6Lm1F8NnPP6KI6arvRrloamN6c
B/z/BJQ+e9yRUxlFzPaXRFUwlHZT1xX65uuqqwVJ8RQA/oiZxdlJe5mHe3vM/PeipEAoHQOCGd2c
zgR3nFUMIjbMfTX5VI9pdoicK/HTzUCLov5GIUDUgH2lrOPpXcvi/w0bg+3eqGWpBqaDFHr5W6ss
plLPTeiBtKwnkK94Yw0fNLp9G8C+0Gk47qDyR4TQIqlxjbKRVGnPvhmzVZyqrA4EgMuAu/YBjggb
VxKJpoyWEUvUFeGJ5goCuhoL3oSs996+FccdLDg4cMMlgSqwqon8oc6dfeO1VLg0XAhwpqwcIUKB
c1EVfmHtMExIWO6NO/xLoVU3Yh21YnStRya8P4ZArCRLl21ut7gqrT/k1K/3l0RkHwQAEOZnUG+j
xsWSwguSq2Jkcvrgl5hj2IUhGbCbDfEhNR8HqAesWnbzUospIfjrYBNOEHVAPWOon2MhjsAD6FxY
dVsE96pDF/gQt8XOkD/qFiawnZ45gTE5SumT1suGyXpPiOVRhdlohYBAO9kLHQZGy2J7fqRN2ZRA
IpDsPgZmGdyRA1RHKDh6VaHnExrdjsVsY5LTxYJHAvXYas1LLwQlQmi9m1S9ClNrTy2JWR5SkLRs
aTMHk5ENdN+eEMT4s/T9AzpnpZoRosOl/VA37QKxGV6/gjBfm2S3L+uuo/WRaoj4ki+DfCdoLSFy
Sf9cJwmkCP7ZmAynaPxR7Xt324itlfuFdlqYiJ1OWgr0vQOBXtzV/eyqaaUJbk/wX6vwTpDnaeTG
eZU6OWTE2zGUuCAqLvASblhH1Fazpu5WMbotD0Q5bpWK7zIbuTyp3L26pIg3IpJ1MQ8TyWdf5BIo
aAz25BP8xOjH1YqdXOlyQuJft3e9VDGhQVHSIMv0j+OGUVLTfTchVZcBXW8nyKFgeRkIn2LQ7XSO
55m35/TWrqhYLB2eBCyvHnzAAYP+bQOyGbXbidTI+geM3gbejCeIAOyGceSMzmQoW12Znat6SJ3m
cgJo459CTlOuB+0kXTpLlDcJKESSioFjjcMAdS9gFvYSTRiAFcmE7kctP3jasHzy9Np3KImIkqmo
D2f8gjsukU9VqYFvgj7BVTIX29SNXrGnXLm7LqiT3UbNsO0i7p5s8jVhofTRQ7iD5YjJf4WhaTQH
k3tip0znPysfu55iFqJ+H+/JnPWboXDtmXGTI89JDe0YRiAm3ZShl8Ub1l2VNmP2Ra+1y+qg2PP8
L7JHqgpiunUwODqQdkiLoFF0iir4OO665tDi3Lktxqc0izAXx0V1xY0WSZCLqeqqmyiSYVdxCwU2
+dDxKHTUSFnWdIQXDV0P66raKppBrfWj2JbgaaFLuV+VbBNlpoe1qrx6AvXirWPCMAIWM8S566dL
3PSxrbxWWSLVXn8Gkft0bIZPnlc+Ge6AlljEQ7hZVHujanVAIpyemwQQkNFc3lke5VmBAMLF1tqL
YRrJKTe2/p1d2GtbKhln+C/7ik7l2OsXP2Zh98kI4Rt111HUlXjq7A97GHzNgCOMS4Hnn5N39o+5
rVbHx8U3r8igZoRlQudUkJ18Oc9KnaWxgqhWYi3Twgsm29+gpb6L+6yBMkUIXomSORn44ptvcx+r
0IfzsCnSAagbv3MIiUbZM3dDchTKzisJhgiANaXmRRk6jwKXMnXhROtJcQlNxBb6cIDcDgS6IUDl
BSlKNWLR0Ajt6sDRB69vGBZu4lC/0ikxSHC6ZQcP1oJJSAxVkuoEbV+1HD8FYA7l+DFKE3cWSuGc
cB65Cs5JRzPTiH9f0CUqVaykwHBxOIRQptkaGI+6aHcv/doLYlgYFC+KpwR0WnBeA6pgvaZGPEf4
CWwTBwmQEKtTEFX5Z9owLLPazMffhAxsxB3Kj3f3noNSsiQFwXW4SlULX64LiO64cRfYbDwwNxKZ
cnB12SviQufr2rcwMeGWM1IGqXaTN5W8+bvNT8QxUDFfiIg05M+qtbyqXWRWclNSbU8amJ7t86CH
Ou+pCgfmIfMQoKT2T59nJaGNjc1/8qjIvOwNIkuX4nDTNEFiChzps3w/FT7GpB666uKFep1NMwvu
dGzRbITODpj+0cnOuk89KequrrBMcd/1BfwCN0n7Py+8AMjTiaRig+5qIQU16udIGvS6uU8xIr0j
cIfSlMkDSymVv/TND/GSbX4/VUEne+2TQBRDG15TdXcYkp0Ym5I8/bQOENRaVlZ2XSCOVWEtFY3n
o+KbOffxKJ8I+ziv7loBKN2lTW8t6YT1GH8RjmzDikh4x1K3pOPDbfw4Duqn1OQwlfd7OU7fWe6y
hen/rDSs3ncvhZiVTtrrWjs41jn9wRdeLJlzP8Kq/2DpXwzlHX38FqKmCEyEBkGoKwekGHT31RGv
KYqNE82qeZi2PD+3zAYqV1kdfUQFK15zvHZfY7w3z7sFYswDTlv0a0aqux5AP8gLRAF+bDPHzD+b
9GZ3gVBpHSiEXb7kCyIgdyIKViSCzJCHwWwmMkVZNNpLgWp74aP8AoibDw2h5Sf77+b+rCP1H/Z9
JXMmWbgWiM/0Y4c+zwSYIt1sDJolldaI8RH70xd3T2ViLdrjJITuJQaa0UGq8sjPCBCgHnOg9lKh
1Zy1WK0iQJLmMrmUoTW+Zimf2DJ9ihb4+8fJ9w7923E+eOpiTi3Ao+oUuK7xl1/7KnVowox2L4KF
EmkIZhEW7ZGdYZNGtWLM+Rky9WsC9m06x3GKcTEIXkcoyBpMrm8lVPQBEqG3CvVtVF5IMNreDgxe
6D6h7sh8dwbntZhAW2+avx4Uz7xz2jSB+VZ412mFV+sBx5CCINiIBA8TB2sdqLNEe1eEO6vtKRqD
gdFNQ5lZ2GCHrMALLOuXploJWKyyiXWi8FsN7/v+4GH9vEj19aCmUrHio+Ch+pjzpZ0EshsJE/nK
vRczA5+qUm16z9YhpnO7UEsqrX95z1MMBHfSQdsDOKGYcWpyQ2IY8e4BgpjF559QO/tfV8Wce+Ld
acJb1eVnEwTa+BpcxaMuGHD2OJFyfUpnOlB/cobQPJWca0UPT0ejMB/x3iJSAKAyvH5SkM4X4O4t
CfS0mqg4TsHeiWmitOjLm8OSDkTkPioMAvn8Ll5yAU3Az2bsS2p2odNmMjyCmauk3TH3FCrI/ls8
dtkIObSuuiNXJX+X/L/gWYzq4gA7j44h98SDutEYbUvUhbsNpPVd7mrU8esXcn5Ke6toCHkJEHYo
Mt+0vFD50tPyuK8h6pnmMKqJwA8CdaUR7OJ1CTVfcAghLgHcb0MmtE1uLrko5nPnBazL7JdL+MFc
UX+/xcF5monRQwMQU73R6MvsRr+dVm5z81/bwN0MTfvCs1mE/OWONyL8il9ImoLH5kbbKSTQMmT/
8VHB0QJwJo3oJWsTmvZELQUSt8A+1+4KGueNNtN/+13JrDigjeUoTjbqs5It04eDwPm22ArnlWPe
oXnoAXjPkE3Oqv+WHcibMmzJd4XMGOBEFQ9hSf87WfshWgfAbZ1WbwHFRh7NJsmTDAPJPJ/Cu9qB
UGX2J4a0DkzvkoUTvjGqxkwmq4gNQGkkgC+n3n57u24Qk2gzteE5oSrz3xzlORyUwRiJBaMABT9F
x/3+QchPDEE96chBO+NKMYcaMz/qJAkcVo6fjYgY0uWL3VdhtImVc0/SusZTh2heFQrF9bFCuOX0
h7I9PWFhcldpgdf+tsYz+Hz+r9xYFD2Q8L5xp1sXP5pvPNLIliPUuHtyZ9nM3ypLEDqppi77rbY6
BNvoY9QeU2gr+1LnYg9vxLUFR+I77KPzxaZeym+rNOHPDQ+7H+2ehIoRHI8ofH0i4g9dji9VjUQv
H8AvBT/jUYKLaWZJGPLappUTFfiSoAG3poNMWQsEp4uOv7DAhbW8G/vCO3uOITLH7GgAH4RVhm23
tVV4AzR0EMUwtofTkLTQYFX8LWOlra8GOtEuQY/hD0QMqtEdGJf/F8JtqHOsPl9pLrKfT27tqUQS
t9pqCt1E9fvqC8Es1QihvrND5PRCDi3QSCTFs7QtOzwYtM703XTofPhvh7km5O662t2eG2tNuGCd
W27V0zNbhzx3a+udkrIpNudBaljZeGUIvBvI4dSQdQHjgh0TSCRmq5K6Mg0cgRHwJ90ULbXfukZF
G6K6O/MAPhcg71tUQHi0q6YURQJdBxDQJ9FK8H4H8vuTmsh6dKlESmrzZMaMlPk7K5Xu2JZ3EbVT
uS/KR6SNwAmc6E0A5EwYZQSCN7w5qRMrRVrVxHMkWkemkIDctddShvwntotFnKZpxGA4M7D/CaF/
cc4qxV96Mvhp0qJzLI/2m7F/TYE1mMeIkFOfid1wTk7qZQ6sD6LPFKzc00OGAw4VwPJO/2e6P02i
F55NiztE2tVfCVGUtcJjrMYLugqrNqUPs2WHaXkYAh+gQGwnpoRwFushWhqKcExabn39lYMyuUO/
ng1W05v11sy/Rp15LWOSbIDh2h5nwyXiNSeKugyOY5I6hpPpbhEku2ToAJ6hlLNeAZ5uM/sOZXna
1mXWwfrTbSlEGqmdUCg7WgqNDkQNdV3ebVow9g1/20TwAaSD4U64LbMxk6QHHpS64jBrHYhiZzf2
4ZlmzM6jxw4JHx+BPJTvSgngGagf+RZsHaV2W2fjkeARDOBhlKdajshAZsGSsM6S9CIUbs+7WeJI
lbnP6aoUxSa/wlLd9OJ2HErnrMvbfz9OgR0X5hZM4AofCFa/6+iY7XSJ8t5EU9P4Ye4OASMXtJZi
mInDVrv863xbYfKs3BBpWLF7yIu8BdNs0mEzAf7pxmj55kfQbSb7EOtSNntDHEcwys2A6znwt4at
KNPl4SPalnTgZ0siwLLvGUypG0Hdq1iAUJGQ2vnr68/OFlPgBCi/vSxW50fANZkYm2mzPSQG6ZhO
VvoqwMdCMXqKrmI+1KE3hlmlU6LjHh9yEda56GPvpJBeUw0zL1vYnsnWUqx48NkpYeFVcEnGpTjT
qwKvs2amVdMGyRM4cmxA5Way7E6tEyhJsUgnShnkWZTYtDAgbUcVFupx+g4oWelsxK8KceR9oeUf
SCiOxh9YoYk7Xy5w7e312fpU4FqpB0YyfKNmFNAWjzfXPTcofnj5vXcDf+vWNPRoqUPmbh1dyyjz
5wG440R0oi7BlILfHIJUVI/9GPZy9sUSHyq9Rq/RcGic1U0vIemicadOhOQUUHfrMmTuTcGtMvA2
Etah/C6iW3AHyCp95pyf2pyzpivDf4VX9/eH4jlYabtcNVnDa1wn7PlVmv94mQs91g6ow7KkT+IX
zl0KgFQIwaKBDYexmDj0tkNU9SEc9aep2EZkJnbVguaV2hYnC+0rwQPbPtljkpMwhfu2hyFQ0cNn
oiX50IOu1Yt1pvTLyNzM/Ip8OEAuGr0LbeeTiLPI+6t8TU6QOYcwzl9HX0iY4tuzAOVmPqohXj2o
ZnNWo9vEL75rNzj/Rt0xvIHvBVGRoEgAaWO3GdAjeKTfrtYikzHDR0J3luFdq3bXkJhJP3pKMiGZ
0hZYQ9dPkQikXOInPUb5qjI/EkfaWn4bVytuv74kKiIx10dk+BSksmdRa3129mewrAhzjAGG18GT
mPyVHV3sIUSdyzCh2x3Td1FDu5poKicwOlkDF9L9HNmc9EaIVNDWtT/gSFZd+hchnvHSQJrzhoBt
nrewYw8UCTAL7oXBM875WI2EbsY370EUpov8BWyaW4LawdNNsZOkjKOfM92VqrFF7h+HmNtgNYhc
XtoQuOzgpd/vAB3xNsQXKUnFxvyA2iYmwWUEsLPuRbo+At552F744MW++NTR3raT0jq7uX76JZzh
a2yTpCJKzoXaOoGBPPR6pSdlhDjz8MRhpGGj6wRhcjKMQYQbM+5NGOc/ZWivc9jKfzlQN4UaDlPQ
RE24GXjTjdncapefR3dFObcaFLJaIM0V3KNwc+Urp3boM3OIS04ztJBKP/GIFolBRaBr3rFJIEAe
tBXX7kyXQYzjugzjpyl7oqaBoWs+g+DYwMU8+SeAGj/yyyX6OBT2oc8em+dEi1XOg74xdu+qzHeO
TJ64ly3Z5ZBttR0f1+10GZT2WMHEAvFY90DNLtQIqo3P1EsrMgYS3RYKwHP9MCHmtzUmuHypuOYB
ZJIm0Jw6v6OeCZ1QrbS9L6rWbCBX/zbwBsG6yGacb7Zk5Iwj81ukqrDD6YyH1jO2kBHQlHHblWyw
C8i4OHNg17q/GLZZd4aN+IzO8DKpUxZbCv9WUsBFAojLeQBhM5T8GVnecbpBHTeLywapU1fXVo3W
nYgFtD49ExfyONLDK4lCjbkfZd/QXByFt0UpIDlBRnkpZboKPxn2U/iqf8/UapvpQ9MwWugUuIxG
Hu7wQpbEKZ8bxRNewJojWEFBETsEp/p3zbFOZenGo0GNGAGoaX1ctOpjrxRshbZA1m6cdtvkF/JJ
SOom70PRIrGcAwV1nv+fqgNlrIByQLkOh/A9Vf/BqQEzs1atGv9WjtpC/wpyBKG81duSFiztLxJB
oufYZTPQRqnEjDmjRzVzP3wVEtVAVgbw01MzMbNsTSR/WaXjm+qREeq/XjOwPm5Oqflz7OteyfWi
XtYY0Xe+tIri4EGrphYMxwlLW6NGdHzwdHZbpY7rHcZRXPFAOIV9KpTOIwXonNn7V2VA4P/LTZgZ
XftVzCDaSJqlWrfIsVg5WdXZxliiMtXer6pX1UAGcjkuB0zin9NKLzYJdqYmky2RUVgEEjKubUQv
a0vvWszrgRPClPIs3NkSfI0lHkAPMcyT6WykBXn0PFaEuWY4osXRJdFBFYpzv+2RTOFZbjo2pU+M
DCVXe53gfHzm7vPrVaCEd+DH2PVh/6L2E4zMb1ede4GuUfXg4QV4NaXp5oRHJd6iw1pBO4jWm2OY
jxHQM4jRZaahDMOlF6HF7800pYOO2A/hFfu/TOvmBYe2VKZYixtBJvXdF/YC13cOXvkmaPxlkYI8
g4CHzCyrxtDg1IokVF9YzdZsbl4i6k0P53mOH7JqELCEw89tCZPpLqHBgsJD6BaxEO8W2aHklkVB
pR/GQl+s2/jDAxlC8snAyoSaeTUOGChauL2RGIEFja0E+q65kWcnnWARxMHF+404omeg05CoYeqA
K7Ht7qtESgUtHBLo5sfRB/B9Ua1W9rKpNNgGua2osfbn88lp2JaRtHHWOPRAcJZeJBhcgmKaN9CY
WDQtOfRXotdUXSlvln+BRaGmgOOX/Aw/kGLV1wJb7XHMF3Di8YvFGLKUiS1hdpm+JbKXe0zqoPXR
/vwsvVNcU3Fb0tqhKlZ8VfAecw5PgEep4D/Lmu9i6raM4JJBx5aQPoRuFtlSFDplePKpjqwlKqrn
g5G5MylA3J9iow1P6+ZJzPQfs2fW7cKtMkwssW0SyhQg9viva/27xiF9nHYB+yrm/T5/eoG+o1IT
UuJ79bb9g39Aad9FmhXrDkAsRVscoK8eWxV59VSQKrHoSjSbwudxJ9BcPhYWpEdcSwbU+8+RTs3w
c2CHWwQytFvqNFjW9bkhnNK2OJpDTUIF4cCtCa8Rh+8ijECkq3RyiC5YjXgQTurzD+KvvsxtWyAw
RWmYjyU0Gver0N9RGWs6duRiQaGjbSENEEbAyZ23YnhkdTWtouOlpxLQHsRqG5m2Rc7vIIIthYiT
qPqM5IaNEQgZ+ijPS9R58KXU9Xhq16Tt3edxhrkpoBUZXwTYBvilyqjbKQLaHNIKPn9KUFVqms2g
eeFyUZ4QuX5qNmBvekWTKQwYIxDohYNsCXzTFHGNW6IR3kNh27wA+ccSU3fkPwfhj3z/2OMaXXtA
tquHundEjrO9gyL/MYBnRNuzqKtjF5DUw6bw/LkY8OeQ6UUer3qBHVdZSvnkcHQ/HTYYx8JKJafG
MhxMsPEkX2mXQhia3DgvsyTgYl5FEIkfre0r5bT+ZZJns0s2ediPph1k+YG1T0lgmI/dt/xG+rvz
fnNEIMgtMEBls3Jft97agzAtVua0tNpV7uticZDAEBspygPoIhdIx4hH0zx1s/gbE0WpDB3UIzC7
HKu7SxpRGQ37tmdJTXeaIFEQoZ5pmjf65QceOT3XjfK95JWbpvYqLTc9dGgiKUL0Vui/HAnoAqmP
O9uG+XT+YETWDvP41vVVag28ZICw+f9rxxXs6C1pQxi8LCzkdx1HDdtgL8Tn7PsHVe1DbE3yXmX/
ZZ++NBirjy+ur+YQx+y4HQw/5pxxd8/fNNTwR0CK6WLcoKGspG84JhBuEKW9ehxqfimN4zpFke96
KxQolMsOuhmZ0ANKUOZLykhzUkPTSmO1QneQBrCGOaUxUomglwp/8kDVcNuUs59No0V1EQqrXzou
gppBdktym4uoIUfHcc4boTiEKoIYz97EPxEQIZ5E6hOl3RgcttN8mIcDaujVKvblzLfJHv6rrq8m
P+3EeTrocuwUC0n7ZJ7QH+88c1+e+EQJfghMfa+jw+yfxGcqyPG6qin/Tu419aJnBCxzRBeEnziA
X+9c4G4ZR30q1r8heVykveOyZFDdzZ91TO6AMdlJz1WcSVOuaQU5Q7+2a1oE6ps+TUXbcEiYMAdZ
awTk/xqxlThtuHGJ0rm3OjgG7Px9x83rOcG/ffWePvQDF6WmJS8qEVBG1+atUitlH5nIeqcz0G30
rYla/jVd104ETsNUH9SZpMsgFX/ZKNNS8XIy8axiExeasJMt/BwzQzQDpKpDZKP9UbiwKmOM/0iG
eqNrn3Uj+JXKZ3ClxWG2E2YJjgcb2lfSV5RcRO5C7gGBrNq++CuZPb45pCYHrKkIjHlFhvrefgLd
ElMxDljcA69IzH/1V9JDCYYdbDRhTbeAjmhf/Qi5IbYIhaWAD0VQPLEpKqkApsDw7/7NuIQKtfPK
ot2eIlcU4KpegdaFFjbwlNzJlofFWDrab1i1PsO++HR0nW8GF9uYMJejOw0LHHrv18ZFhJihv6Gv
I9rSXMG6t2rZzegU9NmMkZdCG9sfSCtvca6uOfALL380JmMSEjfH9KHS9NJ5suVaRnRaB60B821k
VKcb9FJUhzDy26kQt7kePcYa9exaedlFnKTqCl3aen4Su9vIHEQuD/hs8aATV7L3eqpio5ozFT/F
WUwqgB+X2J7agpc6cL6Pdyy6PyypdYb1hmMjusUdDNjzpCmh7Z4CCayDeE35SNsQ5XD3Ji+SROhE
qaNp/U32Ij1E1xxjfor7vlvBm4q8YnpyoKGMs+48i6C4K/Q4FULvqQ4k1BNtt2ZXWpmHekAElMXd
7JUFwq6P8ylDePmUPlmVKOhLb0Q7QR8G3Qwreg4SJlsKYzQ9LUKSoCmG51OBit6f1ebZj2xVXql1
9gXQTvUvL0c/bRZCdXHs9ADosXv0N7uk5ZBMv9Nz7UknTIKRx/nvAIk+Xc4qNmky/t4SQm3YrvOe
UadSTMzJ7WvKR6zBSTq2JXBtRSQXp+GjdnA329Jr8lYUJHpnWnk3XkJ/bm2z9vDAcQvI+kBcJC/p
6hZf8t9WGb2ka+VIU14/hV+Vpzam5T680Zt9itwaDawtdR+AgeTcEfzrOCqlvageeQKI+iza0eyX
Uay5Ju7ZyM7iOBJt/pFIz4KEykqrax2DwWJzq8SRaKpm4ZQRmjXrVbw7gm7Rw7hwYG91fMicmGzh
CUT+e53MHUDqYnKo+qNFwu6Cmqjj7hKGu4K7Bw8psVYSvvY4mydmihs6VcqT/b2eelsVRlNjrXwV
PwQhP9f9J4v/t0ZGmsrxReis0SR2I/m9YO5XSJOdOOkoUTn9c0LO+S0sAEzwEVvuud8wXuqoGmfz
1YYbR4mnh86DL06T1lU5t6w/du66Q6S/SgOfTP84QB5+DaGArdqIzbGpgntMzj+nOlSTe0uCNyEQ
v94NVmch1Fz9bb0K+SXP3aLLaOmTMGFcykevhYMys2gX7jvgNiWCC06rcl9Qi5ga0uKfqhXUGKg0
Z5Zfgx43B45+Jtq3hzAkfKV8yZZDAl214bz63VpzuPimYsto6z2uOHwQxuo+BaA+/Ms5TOYRJveu
f0nlDHffJ7diQnhiki6eivtNtFIFbTbC4lj0unmJUda9roO3xLnAjyeNkGfG/LZ3axD03C44jVF+
/v1bO/OGBplGraVET+rhyY1MsbhuxvNMzvvasTjIqxeloQqhyRWubxD1sxn3ZgN+rLlcLzmOG38U
B4vml5BcxoHRg1AYkwAHzx/IAPJXm+GQ1QO/TC5G6tnCdLimMz5MaHSthB+8WctG0ZlwIN962zCz
67WhvL+Wbj58mBdt3NAiO1G5BzaFSUEpWuqBCmq2YWdDhoySe3mA7Ia5Ev61fq8SOmdiiNNXzoq4
GRI1g0/+T2pmQqKS730iPVwraCZTkV5ArrT1On3fE8KP4TfPsdv5duxgtjhW8sfu0Qi5HNz6tsrn
8Ug/avUvAQBDihd3CqoQveMaBYiqL5Hd6Z4Aw/JJesXv1Den+zMt74Yto4/bWPVrGLfRMJ5T/xfS
7nKbKesVr1UDOFzBHsBklf72zvI1Jt6L3Gn/dtav6RE46gjIYuj6hdimk5WzOPDkWBGaiVTrOZxv
k1mWf6tm0ce/GCivAt2Ca2GvJ6Zk6t6Ud5PpMcZnW3d4sWfF6YVVnlntZeD5L7tCesI9n0lxe9XE
RXoBE75eajC4stC3l3Any2Hw4rDdZJSRM0BIw9b5mABfOHqkkk/jPRF2V7GDEQl8Wx6ilq4s13U0
t2ew+MXxHeiLhEpNPCV3TUQYzEupNcA8JKlL4MlzSh1E9Ki6T2imccjTbRqXLmi93CoopqCwP6KS
4RwbdMHE0qRjQttpsRYg9JCTbDQaAdUqQbWpkPSWvP2NCQ9iykyilBHDCBrx2F8PghIlbcqCfwRW
gkKohqQLAEmycR6geAW8VIzE1KYV5ryUaatH28i81ZoRhRd79NsVdJ6wjqaEApGJ7LO5DQpQBUKK
ER7mIdK33hMX8iihCu4sUrASwWda/CYbl7KDIasuab7KRo+tvO7xz6Bd9Ww8mGqchjqjajkNQRVY
hsWskaLeRdHC6vo2urKMwM83IL/jIYQJI6zeA/SAxM2C3yipA/wUGpyCvxOGyGBMcW2nNtdpjpLy
TJD/ZkJmWz1L0dMMB1/CCsTnUVuSr3lv13Y/acMKZq1yZR21X3ErUjXEI8jU4APavH9Kcz7m8/0c
p1nkj2p7LhBbIzfk0KXav6LU04odY7dJd6Qa98Azd+Qz/kMuF4KqgrB7Q33xZRGQmhacsHd7OUhO
ZM2cOjylDDo87tw6PFpvbCIYSbTZX0eV0xj+HVU5I9P9JWDbwKvn9h0O77qvlbHCKt3q6/v+6Ecq
2ggc9ycyGL4b5eRAAEO0OTqZPEWhhCgUHIpHcd6UH3AMF8qQwqtmauX0y8LSFHNLekseI85SV+rD
Siw5pMBaPhDkJe4YRonX93YhxnH2/u0GxLKI15KZFr4aMoQPGkyWFo0GYlOc6pVJUSUgbL+nVoq/
X2lPKcHDELTEQByG2qzkKAlW0QbBTY1B5wgIV+yxFtjJeQzuDBoYL61bgEWALMlzCrAh3o63rY3q
otXkhJHK0r5ydqOAMPOlgFx476xzO3yepTgVsGdariBzJfbXUEhnfS17bkINPHkR65LwyPA1nDd0
HJGgDoVii4rlKBSMYMjXXWYrqUCtCK0WCxB2UtXaHWVIwSpYcDyi2sCm63JNXaXDz1l/sN3oVtCL
Di1oHBkybNHDm4KAtmL/nuIEGKpc0qlHiVbXSxR29xQxVohW1L20XbBv5dEtaNN8r/6dwstdE/7k
oMGzG0bTUenEoUcY2H9jl7PxmkTaGDwIXx9zuDYisiZHMTivWthDFNabSW3vOJ463V5aqd94hibX
p5zczG9rH+tKKYWqoEkfoCpAKRW1HciyCV5+ynzobBd2GWuBRNIPLzaksAkj0bZ/wprcOqyUTIXY
INKxk7y+A/DoAHvgX4PW4EcFjHfDDfVIRRiMR5+ckjCzyKvAMI817/kRHxvOt/2PRCrCxpr+JBX5
/j+tGVf3+qEr2LpVFrVcEgBPs5+YJl0YV5/adldovHyMnUtn1DHNkUasmV0hvDQ5NPChiDbiRcQ6
Wy3DX4TNPDLPwf07vgN8vu6r3ST4ut2OpmLkxS+Dy60lmGh4+w8JiYckv7qCEoHY/88nyQBJMiFq
zoHFr2I1KP4bBOx9au0YXxhdL8zbTp2SRtJjR48Y4pg+l+olHzpreG2tr3A/dTNoJ+B0ageMf/3i
KdrmVEfjiuZDFDHCHi2Wp+HHc7fbUp6CwKBVNQrXSenk+6qhEGG9AVoL8b72y34kK8K09vlXwpzX
Ma5705Cs7pSkvujvFMmouvObsXTLptdWmBgF0Pnc4/Rds/ODwmuicDWmOaHleHyYWrQpdFws6fZI
uapCyPEOhpDMenpmpTT/lBv8sk9KobOSSajMutCcnqWDYMV1jwx+c4qxdglkYGYvPEcfMwYgH7Gx
q6nAwVUC49DA1/D/PxuBipqwqlBawMIpUKWRQkDHg4OJfUe3tAkSVOfsE8DEAT/Xrc3/zsnMMJ9b
maMtxY0cRUr7TWjjFkDXKpcvhUPeUbdEq/NAGWli5KxxIBe/QXYxpTXo3MEacRxWdXEwPL3dIk1Q
qItlLAYPl+36N+xnfDRHATF4Oom8XlCaNkqwl9qC81sjkUIlOaDmjny8QbG4VaQ7byuoVV+NTyKM
SWbWjF/UfHxRxoP5aOdAoaY92YH5cP/TY0FsMsZ/16ykMCdgpdJljL9SYTdRSgEAL2WqnCRvPd3i
SYFwZJaCy5So7DA0obWB0VZylcvlxcFrNedADVkkqCPITs+hvRBKmdjdncnVAmqAJtsMwF6XwVoK
bXEywk0cO3JJna6k46e8vKsinaxpH+jGhashJ1wRBFOh4a7p8ZphqtxhW+X2DcXZiHmPlQUCnbiq
n4SRFyHjTkn1e9zuL59C5KT0tk4HsLyMQ4UkYf9v/btrnDRr6wvNo1o4LE8dU02aMibvjbxhdst8
q6wwfI+89bHlkFIoQDX17xxV1yfYrUYHN2qUdcsuYSQdExcpJKr2yZ6VQEFTz+e5GU2EV6a0UF8K
dzpEjumr1hf7k3GQyDEf2EY7ypUlx2YSwDtHAnw6Qh/9wcR5Xlr+5BFT9YQo20c6LTKgd42dlQMk
8S/qoXWI+dmrtj4fWA2IRHlqF6NnXe0klwgHSptLgrbsntt47jfc8GGL1W3b0oJ8ink5g87pnJoI
o2P/63Kr/l4YJM5+S8gYashxuHR8yID2/PEAinXsXghFzbX+iJ+gt9W+PSqUT4nHceou+pDD4Egq
YvBmbXGWZf/BR5z5aGIyTcbmYe1Ko57+hWlr/N+cCqI2/UPj6HURDuf2+RdXHDdwQAVS3jDK1sco
6YxZzxCHs+QHmovzyx8VeHuaLN2qyyPvqrQYzxg+fZc9s5kTzejW2xyZHkOc+J/ww5R0dAbqRQhZ
U5i7p3w1oKULYTrsbh3em1e+0t0fHmc5HLBldSf/GArNQORtYlARgVLjSV5/vabftXHltwP5NV4M
2OREMGUUIuAx2JUKrcbbUyy8nrDFZAyvEPEQ6aAcb8i9Jj56ameVmjgEL1Q1FjuchPYmjbAYragh
uO/UyF69C9wH2zxNSH4IsZBohsVA9GkdK1uRoP5TQGkRwuY2p9UzdfZQsdrv3QGO99RuPWuSHa9e
L+p2W0h7JJ8V6GhOYLczAItXZfR4/jSWiMiE4oc3KlpfuKY65BtMRYVR6VXoGgL+IzmsbwTmDeI+
9droXeOqITwJbtyTyp637rXuUhVFASr8/o7lpTiBfpwCrNa0mHhdvkeGGrbraptTM5kREUr/GlWG
sZEYNA0PwAo5K0bEJfU0BMl4XzM44uHDg7ax5awHvIKDRpLXsCuoTodWXenj7Lx7/omvZ/q1qv4n
gWwqeh5VVlSzWOE1Xi09runofYy+1sj8YQRf62wDFTv/3g899x8ENNDZEqqRTaEZRSkBts9m/pdM
8o3v7KElMFzUANI22DzQcd3cX1m4h8WK5TLWaOU1SEX+9OD+oMPNYIzNaFnNDe8/aaa8EuxzzrQw
cgaZGpUKLrgl5wi3IUk6MNZaFqCTTDDa3JaKzad3mAt580c/ppD6lC7imST4V04ELbYy4FaboGMz
pSIzl4qiSTMVQKtNkHXi5CAUYrRcriRtofMIvq7QkNJI0OCr3wMGiz58V0vbUhA7+qOwlClqLqLI
8BGG3li1+bEiFRhtH94YgtRAE+Hm1w3jX+3kgbfJv0K59e2LT2bQBqQKd8XfAQ3LCqVGfsoXjHeB
Q6tGYkf7YxkzYvIadHUMnGwJEbldhncsyLYd7+t1w9kWIgxKnwvdrN1c3hptF5fNTosl4YLszKHr
AdOSu4WGTjXWFH1Z/GquKYE86+j/nWbEGlbOQdqjaPrX3aZtKmOPham5dpShFd5/jU6FqkHdOfAB
rs3YP82RLHb3WVW0ssnWYjSlFld7fbTmjc6Jva2I5LuNDbrH81n6mjCi5Tlhvd58X9VqoA2IREzE
/YnHSFtRtSiToDxIni0Zyqgjk+0F0vIvpmeLwnne8BCCzm7ZGORjOni8/uaQUQCwfEHSmU4fEJXA
+kQ2JS2EvHTh8lyH7PybQeKOHi/l4X/dcJTvZR8IgdondCU7wauhAxRrh0r6FpdKT26USlYTlqkO
FVBGZnMuwA7XgcXhkw2qXYnz3Ue4i9UNZMtL0SFCJpVN/K5BMfDy8UrN6/+fo9hZySsF01EVvjjp
p4WaobIn2PxQq0rJCjS21jLBKUs86JdbnYUYopwkr/Y5cCaMy95gTBiODsmBCcXhHlTeufu7Slox
d3OH8hiDL7Gw4LeBiXCIAW/kbhBxkXhUh6jJP+bQJBIxAtQuu1AK5EV64/bH+mYe/P4zub0wzq1P
KcxrsTReC09UUxCA36kyN5rVeOQfzQQ+Wpsk+P7CSVue/IeAKZfCRQxR+NbawQcsIAcydDWLVbNs
tINLerAanJzpz0xGtEWexYHQKET/F1+nu10gwQib+1M0UYWU4/D5Ov0U5+KDaT0ENDRWWgMCCdHR
5ukTDh5yyBnFdjpQbFTATxpm1XmfE6AfPbJ/UqvxLLdsmsuD+Rnjw9OVttMxrOfa817UsfyVeZ2L
hoh6L0oouxnRoOZKrphPk40OOrs9g6VvgmLlJmggeF55B6VX3JkAEFZ6aFBR1viKh5G/4ayqBUyb
0kqm0QR9gqr5umeM1r2mCgHSizGeIEi7XTpTFTigz7hfv0goZpwTtub7P6Ko+aCtIa7qZfwmS+gi
z8fqN9Hdw3psXITafNDyoh52kyFcQ8TqA2JnCqG22g0PXxY1aNYvfyOY+L2mjJOm6VhXgmDTDU/O
aqhZn6u17ZWVNH+GQCyV1Zi1b2yhH3Gt4II+uqrl3XYhmH6QC2DCBK0RU7/6lwrhnsNsmpUiDQO8
tlaxNCebDQV2Rce4DhT4jC6C8QIb11YSsj3UTh2ZEEogvSVdTCbwA1PqjBQ1jxrA/JL0fJUnNyb2
yIr2eCWY/ACbuoDiqpnAWZ58Vm9Gb/ijz/T/JxmqMAnVeX5kl1duf/yfqk3/hkf/qqTSItZEU2no
abYG/aGTymU32E5pBMwi4QtOCbeN4lTCQNlFlJFZOc9DbWNgPsQ4gRpoGmmgvBiq8ieF5deGMnWf
mCwYZgajtWZe6GLs11Q8b+j/Ean4suWF3ARW4kbUU5wy5YwI5jw32ObmDdwyHg/0q7Uo1H/0SG/C
2aM4444XcVfgXcMzpFK9lxkwZfs89gSoj859vi3Wc05WxWyPe8ddfNH+qTrzDVdqxqatB1NETc9v
PpfzoI7UiEeQi3j/4xxZJqer7CwgeRT6JQHWKvJuYu+8aaKCS29k5vDvaMjreaturrzmiosOuRhq
cRg3UcdMhK1dq7M5/ZqVxt7M65yqEV1frP6ggvhRmjhBI7Bd0nDMW7p9kA5aMkSt5os00G0IWMEM
cugAqOJjxWnotvy0z/h/guMGiWJmP6XPxR2MRs9PPW5vjfKIh16aOSJjo4/jxOQChzgLJ/FczCPK
m+c7yXVIlUXpLwD5gJEz32L+Bx3HEZ15I+wqvGFSCjbsuk6sVc4UnTdc9Nt/XmqkC5GwTWkrha6S
XaxwuZMp/AIgFDBQMI+8O/XCY2WCwUfeAQELX10mxfaBNZqLZy8UaZyO4UR90/hm2CedMD4siBRA
7YLr2ygy8acc4WhEE9WsSKitZ38Ipl0QnR3Qsyjsa9kcVvGverQ3b/QvqSDG3fiaciokqhL0LY4K
tZCyzlMuG8sXETZ/QylG8LDwZ+MZgubuMRY8unSRzB7cZRIU2qqOq8UcHpeuAPEVIr8ISLIGnYo9
iwxW2GsyeE8D4trw2x7DLymy8BymhTaC9wCbwW8V1pakUaVZ+N9dzILnyQPnajJ81pW+0puU8ctg
rjbwzo/PwR2KuZz+MqfGwBAkdG/tnJkVh9Yp7Bgmg7QAH5+TetWcLCBxSSHL3MEypXYOMKObiIog
10sXUTy/lfd/TfBFEzqE04/hGNU1kClBW/odx/gw1V+2ePGX9ceymLn1B4u7aTcFH0VskHqhMTE1
9H+8g13ixKulU8zTMLwietptQIfhhUqXovcFaTyrwDSAyBfpocmajCoHMpdUbNg8ii3KegMNdPP6
sQPRqKeKpwQ56NAny7ZRr1B31ZFLnFUgvvUdaJO8mg+KatkAHvPw93BIciWyhWPFn37Sbn6IyXX8
AzDieusCxABkuVw+p91hsd+29OOVk8usTkFSwOqjVVMJ2YMBgvWgsQno4Z/R4KGdxVZAeE2bRvs+
JdpbZwY9gKVuu1La1yxz98WtnSkeV9G88GJs9C7okMBoIWufjUDcUCjIHCy3B0AdLFNfp7P0hAyG
zbHp+MrhCFiOZ1t+lHMhkJvzg9U++DEuL4mdTUndesHeqosjBPxLPkwNE3p1mOyag5sxUlXfYUDE
rrrRi3/EebDAxVunMKhMe6kC7LwxXQaS9AarHZX0xxJ38BoZamsx4of/V36gjo32rszH3IWH+1hP
e/NJdrhzs4s/TczsFe6dXMyiaz3PxOmfCUVULAdTgckGlPoo13bATn5n+3CjU3AWJhk+ibohlF7m
Yyf3xtlgzA2unkWl9td436oLWZWqRLfvSGhxbnmSMHdiKAreF97QxahtUfbXX/nYhJ1ASwQsJoUT
vBcyFx2jhXsuL5P41qfg/x/MbdAZ1DtGL6LsUD0TUGkt4nh/1wCZjyLTM0iS4dUwYCs8WQjeSyKa
BGhw3J6X8WJXM2VUgHNwa0gC/lGX/UZYg592Y2RywCLn24glpSKwQ7WoO4Ss1Y+7GUPkH9lEudeX
OgmYj3ipfwrLh8zKhx4DMlttbJ2vubeycLG7yASuAApKJKCpaDka3F/guRn2qfx/SVjbLxzr3Vsh
HnSYoSp8VIH8DhVArYbdVpCiuY2jWd57rWDGyDEYVZNkqD1rYcMKt6AHjUY2E6TcM87H+5HCv9xg
ef0m41BvhqGP/HlImDWeIatPrTqLTiBNY3759fMR5QMHw9z6bY564AD7aBdWZNJiz9cGSPpW6p8R
1BWO6S5FPpPNqqY5lqjmOV61AFJCtkgtZwcMXaMpUTu48pzBXI7ex5WlMLMI+QMd3Jhkx72FRskK
riua60ifWRJiU7435WTgwIRpxoglT2Kn5LHhn4elIZTRZDsmY1W/QrPLXFtAIyNbUf8XA6dDd+Vb
JXvLuRIcUNE6ng44LPKLVuFh1oMBjEubHi6VHHd+FAk8wFtmQZQ3sgChdBAv2BkSdoR8FYZTFGWa
HTWJqcPFmZvS2kwKJYLpASvDilr7p5Fdnhvme/PiJmM/ncsyDdErEy75oqeFjM0km8sTyGBaqd10
CrVuCVCjJ5xpWgoExFPGaw+b9SHfAZ1egTxpNm8Io4pt2CtH02nj6IFl6F3aUKscgePqs6cG/OJz
GgHDPJI1kkycD/fgpTi2KF5o3jXCPHzoYKH2Ve08KFCzy/zgD2XNQZvpfbiUyPRJqNPzLFF6rNVQ
b8p6+dZ5+925LJ31KcVH/2bE+Tb0iTbGz8bWBrueQl2SQwG3/nRonjiTci+TU6nYUQcspBIot0of
gfeW0ruP7kGxQ8H+oKcw5eaYTg05z2YfhSw4YO3K8H+xhS+IRkXiOos7OeOLfFcSbG7Bg0QKheBY
DMKx0XHjdmutXVy94e11dQ6uPn5ZPqUv3VL6h1lAyZSztUlnzM6ZlipO6bKONIO8nSCvMoXEJ5yj
6nINGlYKhAdGcbX1NQhs33rdY1D4/SHM1QlTL6qvaOp044Og7STiEE4AgdKku7Mx8BqaLBwiFYiD
UnAB5+K5Qfiz8O34+IkTPdnFr1Oq5sO2JiuyVnTpXfu6AKpbZOk/woRMjAjOYPGcmjxIVm+5hYX5
ZJCeCIwq8PRDtKelbFDFjYoxU4YRKD1gaikQnae7aH8xDo8WINWC8XZcza/jy9OqD7wVE8ZxG4FL
pI5vYC7VEU6GLS2HZniyOPmldVxKUVPig//7tdYwgGfyOe7kZYyZGHH+fBKHNAuFVRCPVdeub4Ok
4AVY8XXa56wu4ZeGAkPaX5DKQMofbRznZNSFR+A20aAHoHA6+uJWJr6UuqNkorzVCUDHrCxq4xxq
6Qr+J2dzCAOYPAHLT/wdvgJVrrh4f42d2CBIJCe8ulsH4SMvvSRaDcXne4UCzKpYZgZLCw4YrTga
jb/qW03cmKagk8e2UvnskY+W1riz4FoXxChLEqMWEPEEkofdO7l8UOhTXUh71vK/MgPtvPnrkh1M
S7R+iZlSjWNmz8oenlsL7aWbyB4cVeDIJR0BGn76HuqdyHBsK0Qks85tNv/Hip3f2OoFa+NBCDvy
TOjdDur0lbpIHXfCGyCTXsHZT5m7MjNx9isWhdMVAyS9DP/9AS+bm0rqnczuLHOmERlkuhKFPuk3
K7N4IQX1VH1KIEkD3i7ypsqZsAGDmv9CUoKZhc37b8Xe+R82N1gzm+aQZYn5ZHFpvcOueZZG4DGm
N9uZSQIcEHIjVbPB+KVBkf0wQBdoBhWTwsWfKzB7bjUaOhc+D6RyTy50ftsehjsTpy5PK+kbVuf2
X8RJHt+hsaJ2jR+SO65cN9x81LZ0L3wJECTULIgiMsIMN+oX5QjF1MCeynyyCXsj878udKMGzYop
BqtPgVRQOgg3ivcKozbDgJOU3tHNnzF6eU8RjbdHFpU9wghqFuM0EVzBW0topr+lmrorzZ2ZHCP2
XkjZthjmX3kv6WOkE6ELXpYuIgcmQi+bovr54uIYBEH62+0oqUxEkk+wznnKq5UN891hQ80b7iYh
uGBhKFRO/w0Xn6beGXIFruSDmXRGkEyIyeol8DT0uUpXvpLZVLJJZvVIRH3sDAUyBgezMsF0RuCC
EJ9qnFYYJd9nvTXcLJSSfgrvflk7B4zDyRmHnzntzuGeoZJTHrU/f0Sf8JSRau/O09j93/1E1YSg
hJMx2AQtVgwd5gJ5M3Tp5nu5o0YDGNG/FZ/ON5/CSFOtQ8xX6hiN+byygUQWiFKKhKNpjL6dlamP
7uJj1/4MJ8Cv6+95WIFtLLg5wSrAn3iAzpgfy/nAuNKpoP/44JyB/9FhftPECucofJLTi69EW4Fd
2IYT5XftEcSJh0ZYB38szYrO705w1x3Aji7hikjkWu60jwvE2Bic7U938M+lT+CEryASFsVYecws
Z/5UBorBrm0XDJYDvltoHbI2Xan/qos79tjQSb5VLKgZRgPrGd5+E47vzxWKilhQAi2n7iYTCIlZ
r/8E7SfNZdFQIv8Wwi/LiA/WqT2+ZTttb6cC1cnIA0KQbkrFN+P3o8+fUpOKzUoGoib/TXxVOoCj
a77k+MqgjDlQAxogo0MsVdo/5bhbQxlI/m6yu5kev7d51IMamUC9pNU77Zs7HlUnUWkh5el7WQR9
IFH5J+m23sHAFy5mYaQJENZy8N79MZCEVYH6iqyWGT5Ifxmv29qnx+rvq1kBc9DXIQw+Hp4DC/Pf
900wkLommQ/l9OrGA+K9elywWCz9eWeNjuHW7wg0ZXYYTxOrQFk5PxZu8nMEKW0OqkU/KLFQVXD3
ejENXTSN9yG7KDoHMJxyDFWyH48uvapwus1VTF5Ybse1hlwNBIDSfQ5V0SlcEMQBUIANGMkpsgzI
apqB0X3Sn4no3fNcO0fyiv8GIjdkVfNYaBkYnPjc1VK7zoVSodFkC5XnD4kYrq4m9gbUBiRkbj16
oe6KrYoQ90mk4DO19As45Quu0+lPV1RVSKSILRduZqDeQUrhoNoEE0Y6S8j+r+Wt2UtpSUVrnQAy
ETPqVAwjy8eevlndB/pj46ZSnOFdTcvK/AoURg/NPgsrqonuWW4XwcjXBLlBJCvdRcIhdzZ7oL7d
mHZ7A5nubar06PDPdMWvY7MDN05SvkvTXbA9x+sx+re6KCKwcFutoA9D518YK5JvteFK/tzQpTCm
z65qSqp3W9ayFBSCNu7p1G2oPm2fU565iQ8H8hVl74EaakAlVBQ1a5oi9vMJXkTcRJ889uScoaRM
UwiX/pTYUoO/lz1N41+TA3DrB79fnzWJWY9pcRrJ2+Pn9zbDleupOTQsocH4Qt2QmVEE8fnuJCmj
zjq5WMJVVCX48O+q72qdFFOhOOikfhCh6OeDskN9wpCaUggPA5VxMFDBYKdKAAosSvckrTj/5/PL
tM1ngTiWc+V/q3tHGilL7taWVizPIU6HnbZUn71HCNsSOdwIebdUwfN5AHtRGgwIL51CsJUP707d
u/B9Qm2c/UpBoprWwTS7+xAK2XTNx9h6FdgfZ2v2wIBNAus0PJGir3A8VeKns5KwBBAUKg+13vrD
p/g1epu48cBvDd0lJiLLQ645Fu63FPLy+Xw27PC51bl2lGrsgfjC0OJ0bOiRPT4hPQabPd9YID/6
KeMPXTONThHDEnfANyoErt02zBIu+rqc3QSGjkIaDgxGjiZ9QOOVnd9SHcS73QxdO7gxHR/VqHsH
Kepj64uaWqMLu+Ll8IIv+EWFEi+mczHURMeoJiFi2709vqMbqRNgWJrAmRsNm0ffcDJpFLYV6ukW
8xv86PwG7nBJCYv9euGsHo84YQDB1eFIxBiJD17AWz6yV6z+KdJT3EUbmSAkSue6BuD8NrlGQbge
f+b/5sKqqEQBXoL6UPCuuSvqCgoQVmTvuSan1QsCrTtu4ztUqHueVI0X+ZrALwvSSwdqLHuywk0P
tiGloHXNmdYOFjZOE7Zhcz0C5lxlwT7vQBTJRWASUO+CMwhxSU0GPaiCwFMhLpw6Y1ilDjB5f5B8
TlCz2M4WTB3gmf1xR5elJYkZVicDmmCs4kHXlNRHO4tZR202ttan5PjzXT08Ee0w3BFshzdMZV0w
jLn1aXnqKf2IcbgDwoGm6xNe0M3hiblu/cmgxw5OBWEhSgxdieIs/12dfJNzjKrwQzWPxaaVVNOx
tS5KzlBtuz2BKEUB5/jAxrHFCsgm/AnKd/2vYCmiNSfg/8Cfvk7AGj/C2V3yqj9KWMNPvcLmxPYS
9lJKTsk+Z7RVGFVCDZ5PV1plrmUSjOFoI3Gnk2bG+V+VpaSeoCi3S3eyGc75kaRVlsJx2+/EHdzG
VVaVPmo7VrISI8kWnp2BI0APFPwLL22RvDhMWA69fUEDH2r7WywgCXlqJayslubrtJo5Ro1fTyFH
48XCkpwFtDkKe70Cl/qxsewI/M7jdbbWbdQKT2ONd2HD6a4kx7UtqyYEQLsC8xm7gQXkoTup7Z1i
lMaZ5KcKB0dGNtnOXybJZW6y34VEVRmT6hhA+vjVtRACvDjPgqxMkg+rl1XQiRvwPfUzQOodtLiu
C7YpjIvYSAzn+DngcWOAx2iJ6+ENfSFqibmDjz5LeTzSZ3BmrlB4b5kOoKRjuAaCVawkNpkTm0CN
t/A6vLLYo4KLRfL/kDeQIm0DvhkcZAkHy12lXCXGwMOmMAdQAX/isxpGXBqgSR44qSyfHzdCL8NE
tJYho507JrLgaCo1FY4CPAa11KWYokTZFCjyRVaot1YejE348E4K8yebCs4nGaM1DdcCSnCV/oVt
CQpEjtjencxRNbHUfm1vwKldNT7J2l/z2VqMvgQjJsryMi5LoqcLnsRH2GDxvHVclMjzZjSdclng
jiOg/R3iyIJLRNJIeYKIIt5qjuJbEO/TUwdhrtH5quSYVvPUff6oZCEdj96D7tjIeepsOeLgCNHL
2A0mEz7oF8KowukwpckdAVByfgSIVAqB0cFpgJOhKmnj+RAZxHivuqmJZ7SOOtXN0Bcu1k7QCm6X
N3CdKH5/YEay1QdL9ktxyjwaiOg1YdLG64dHOTLTZu8ve9WmJ7yNMpovQAkbL5+MRlSDoomGX7aJ
xpt2wv7PVSp59JQOmzf7maRGSlGvh/E321Wwu0iz39GmlQ7TmFdkIxuhI/N9tZDL5v7SJ4Ff9FWl
WBGFbc7r42YMmOnfi/lt7+ouFglur4cWMsRWQy1rXCeKZCdpRj/Og3k74cQLp1jwimSO63gdoiKV
82/TdQRH8Cb1O9i5w2Dn5exQs84ekIwKasorlrKeNqJmXyFgumnhm6/DAhgU3f2uss8O4ykTJCql
BnkxK8/T84BiEBCGWfYyp9+vnf661ot7L3BL3mVwg3cZrU1hzu6XEd5bUiXWsIFb1gBTGzHsYMKb
jYd8AFUwRMwgSQGwnigbbpjGJ1zOCOEHAU2auBMxQxI2cMR0hhSz2S1R3Fw14KL8f0dq6ZBxxYAq
9QxRhKZuD32biRH/4+sYDzW8CSkoYVl5QBoZ7+015STaKhZj7QNJj3J2MBQMloRnSss6ej0INNGU
FIgHO2XXbococyiTHHyp491Gf1s1fbLN0Y8KZbROouYiRPydDEbLKxLywkVuwRDBa1yseNJM9dLD
uwWRgDDwsFZ6bx7N8O4OTfms/CJYVCHC5G1h/GV2BXDxOnmRZduY0lXLYcgCFJGkkieFL8bBuXJc
t/v+d2LK0WKsNig38aKd2tCUf0CpoDC7dBkJ4Vxqs0O+hMPLqtvbx2dAepK3MlL8UuPpLtZdRWz2
6+JoCCuz1+KXvY6HDrSczIOzMEv9txNaxV2ggOJL2GNaaXRewY5WICvHsdiLqWsTcmcMPrxuGmTH
/KTKsnIbeQ8MQZv4GCX3DhQSkHL7bR6DxUvR4fycS8kpt28NWY4dA4gh0Trb1dm3SDnHhlSPAqdg
Fd74phw0NywSwtzyKVddCrNSeRQItEb9BCu2mzEwB3vUiprE05lv7ojSEulNC9za7IY/Jt4d1O/t
OCzsyMUWIMK+41/p4XQ0Xmy1Ldr4bJs4oUY2rrER1hyXX24kqkSt6YsDwYdOviSyBQxUVe5ZsgZ6
KiexGPgNKAIzdPRBCvrpdTqv6ogO5TdGNux79C40ljhhhlbLRNNSSSIigsIDS79J+flIBELKake2
mor/4ausBlok0vsmsG1ZOX0F5DHo6suiOVkaIkqYG53NSHrZmBWcUPiabXoJ5Nh99ZfLTbTbr+rl
kDkVF2flXtG3LgTJlYMNUPauTqEokqp4Bh+fR6BtumDbDnsPLG90115qEK5kERdAlQuBEpWbSFqa
RHTbGV1JjJJiDxJVnL6I8I84IFgQFA5430GG/qXoXKBB52nvVqP4/659v1h7dt0JHIuihJkmiUah
pIPrJGZyrcp6Nk3DbA1e7ScoINnOTL7HNmyGwi5rrVLECwNUlB8QtJjW6uunSxA8rOf0JNlNlgDG
0iX+Lg3DjHFteNhbwzw92JfH6NGP+K7Rjs/9zVgA/7cB3FuNjO9cUwWPkpLYEWbF8LqCzyQKI6g2
CoLPoi/yFWlLpZ6asL8iPNM2g5TGpIGUqAv9XW9uXov7KLwkUM8toxmzhIfqhaxDbdZ1gFqPuGnI
O0SMSoVY6l3oZ3UUTu41mSoGy/XEyUkxSCTXF/qTmfnBJxrXVPpL0mSG48qnZ1btlvopXPWzxlNx
OBYka8JmmvQv3kQXKHH9GOCnyPhYTujD9ogFKKqngN1bKixbhtHHG3b0bStj845Vo0UR1oMsgLbf
EZdTaqyVCSyZeBBUqLcAVHKDABOmGKdofjKATqz6J3SQxz+cwFsqH6ahdqYy/C/+OniE6GhZVZM6
duG2PYkYTBmUkAUGOpgX/xCNBgAKylfbIQyV7SE9tKk9RWg/+0frVB00AWhNLZxRDxuf+bIh4m5g
JTczeiGAh1uGXgP6+P0nQrBP8fho4oEHuflatyewyY0oF3wb59wqcveLmw9YAUaY2Hnc+ASTShoX
GEA6dZiPXjmZqquU1o/iqsslxfz8G8Y0Dul1QCr1Ke6mf8rP20WgfSZ7QAPXci/4N7jzJ5Wz0EDN
uQx/UaQyhwvWSYrMpDsAL5K3waUfBZaO2o19nDSXpp7N/k7LH9YNfninOpv1eu3SFjm8cDxgKCm5
T+3huBFxDNPqoX1zVCfpb+MbHikRwGWBQ98ui1afcm9VxoPqLNX/UuvxdhsUBcljVShI7uQphVJF
DcgGfIUoDCR3+iqB9Azdexx0gaXluanxbGBwh2PW3f//mJa+ifuZCdnx+/CiRkGUJgQuzjMH6Z7m
+XsW49MdiCJocmxgeFW1xU9IA6X77n4PwHI6ubNsUFREw/ccq7l7KPsY8OF/kaxxaNGNBz8VeccP
zb7Cb7lneGn/ZIKJZ6swAFTE+QqLr7+LlHHEoKOobkSxDKO6kzwyDd/YROPJQ6qPdxfsqBOZIWU4
deYTkAlqyYCxE1swvi+UAuL2ufnXzaZ3eX8KIIUnjOdmRlvrRQKXXAC9Qt3JjGD9/Lvykoip9J1N
3DCAAirs3ygM3WtnG/O0PSjPfzoek/nL8WPNxSrApLlPvLdq6uXhVY80Iws9UjKE/Yn5yCkJL+Zj
2VDN9YSWdB2gjAwYTrKSN1501p/u1FvM1wm8jiOxvSRo1bJz28+TlTdNnZChl/VKMNvtTys5+qlp
HXeGxzYdpcB/2wIVjiZqOFaiuNyk2fBuOqnmLgju8hkp4vqXKBbxKtcB6OHrhx5gtjhpuG4NaPkB
HFNi+ClnZpGlRj+xif6/a5Ex285u6KKqyvAnIMgfZ/sx8Xv+w+Jp0y6lMsFL7+yQAlc3x2S5H/J7
9ppQsjvYOdIICbvuZ0nasPBgR2dI5S0JQG3fb4LnFNA5VSjtPAvCx0fusaZUiJI1LqPfSe++yPea
szzNpOxThOs2YkaHIUS+OwEZ792yqJEK8G75hs8TrJuUPbCElsZRNnh2XSTaU68tciRVKXdEN9Kd
NgG0K4SO4NlrcFF65p8SmIqdci+bqGphNaq02IncEC5AqK3jSEgzSBQzQTS8rPak3Il2iE4JbYiR
SmmBZccjePc7CnJCUyQ4BdG+pw0lk8/798+bbgnSIUnz7R/6oFfgWS47ATd92MVi2g/xt+mdL2NW
U7nlBzj0KQ7AtfZiHqWqN1MRCyaQtmimXiXDLW5nHp4C8C5rI0tJ7cW6h6tacEebTGsB8dhW4yE8
MG6zDStIJxPVCurwPqjyCDhll2jGS4HIZtWT2Q6sG4Ja+aZVuGHcIk1y6sAVeYujiRXrHyGbHfaN
t+c3OE5lvYG5OXbbe5arvd/kkg3CDPWtS39Oys+xi3xMnHSZUkSqOEbiZwYmqH5yWcxTN7PHDVkX
Mbww4w72PYTsvMD6gWZm6CzliEXKDO0oyh+kvUTnjxbiQAopgfA+HsDhgrhnFPHfOTINEKxjk7Cx
mTUy6I6VhaNsU9NKoJrEhJQTeYfT8GVACbNFBVVKgZhRh8eHMCWvZdAhSn01AME7sVaop39bR7eb
ldfoB9MtxlKdsDE3/Y/w0IjnI4X0F33YQPSmPNk8lNlCI/PNFaOD2DAsmMiHdqDEJIj1SvcPrshD
ZHdyAsLjcLSy4i7iyJT49x4EF8Dl3x9AMK3/KzLfLmUtbx8MsSdZiChg3ejXeeSQMAziFBJ2Klpv
t1qy7hg1mf+sCyFWt+0Ra5VsUkMWCSU7Lr/vW3YC5wkb3whUuXqihTRk8f2ZKZU9TElluiBrw016
kpaGsBm6evtF8pv90/JfiGCCqGMEoNiHvo52LwfTxM4ZLUTSJ5YL3snXIaQ8YVuQTxqtxncsgpgj
kc0S3RrBFextGCSH3nzeEiLsF2TnQT0lf7X8cBDLr5vIgjxODdWVreVMXM4oFzXezKIj43Uhb0uy
V3V5b1PLQKarp6jsIMjQfPmvWNmdL1lQ/UBRuv5ifb3JhQwli4s9W2rs8jGJXROoHuLZfIoGXIvS
aHICN6OkHuDz0ESGHOZL0sw+dkjZKv1nPk7Q5GrUwPm+v2jafUWgL6iTYE9QGRPPsLPncixiEtnK
B/1x7YaIdBjOFbhqobsM9eFuFxWoERMvtDa2HKVwgp6lujm2KiyvDoK3YNJK4jnYHk9U7ylhpfMZ
uSdCQOSo4jUICKdoR5VG1FI8EOwCLK1JZ5MWb2e5OJ2SxZlVe3hC9R97k9csKNWUAQXi6GucJXcs
pCPdHaYWF+Cyx1GMMvODgfOYf/4Zd+ykuJrK/m7Leyj+15Fbb41WSWLxhWJRvRlS00MHMyPJXb5e
/SjesWnY9/5ldV3n9LfKAFgKZmCephWmtPs5oE6qDM4MFDBmgBHv9uwRLzFNhj5kYB3wXUQAs92Q
ynJ4f4b2P7fJUq5O/enh7NTJn72Sc8TbybfkJPGgyPO1RX0PU0jx9Q1o5JEip9TxKzXRu4uxmVXJ
W88ANC7bu2sEyx7gsiD635gaqwDQw2KiqTdu6CDzMy3OPp41YSeftI6d/fhVVWcediI7DF2ZYugD
8uoTcJUxdYnHDgZm39k01AA/iTjaqXTde11pGPlVD8WtYllWD5Bv1G7HKVFXaX3aaS8EyFcSzPzM
CwSiuJW1/iJkbdf9j1rvJGz7AdE7i9xjqFH+orO0gys7K/7mGe4W53+GA3h6yUwoPQlDo+1V7Tt9
WYezzo87XxNYFheleIQQOATMn3XALcYPotYj+KRSMCC0XjWYtFb1KZtuP60Zuzp5na+DH348uZjl
481rTK565I3lxl67TlEu/m6Bg0yEnTXYK16l8EnL3a9ilvILJfiVO2vv/6pgLHxfXQTrBDe2t4EH
5W5WE2BXl1GSnlVf+GIom2+TrY5mfJkbuarSqHdIz6U+sOu8k9DtSsP+4y2Vih00I8i5kRiSSmo+
D/e3vEgGgeBFEnCmvSRiAW5nms7A1zDX7x3+940KeN7tabhS3hnAWBmXkjaavH2WwpYEwJQGJKaB
lCmFprl8i+9xHVvcQokWXosTiV1xL7FCyGyfMAMMgaPqgpwNz41igOdZjA7ECbLYVUaBngM/nHWV
+/JKozILFxBrYOGqUpJyzw3sbuT7rKMzMf4Dn1VfM5JzmCC+2/egZWQO9qRTBX1cF2riikEPbXqi
U5h70Ul6hMk4Z2mC82mk5PUezKaHljqDNrOXrhbSvk/o9sAx4fB9bVS2wg0+5rvWm37GgBsED20N
CsNrjP81MTVU3Uo/1i0JtPPEj4BQkoNN84t5Or5PtugOQ2bNqUJk6qxFC89EYQp4WraUJA7y74aP
mNFtQjYYH1uqqP3DJqBh/iDYcGJaZi6D2G2nYKgEW+OjYg7q9Ujm/J8tCYJ7t4EXMT0w672oQQcv
xl1briwdSdyZP+ekihX4BfZFVJs0u5mAj3M5E0on3H2DxGCGip6cRFaS3TV5ZCZ7JF3Rybrtjzrl
2mQDszk1gXoZpJNWFjOoRZlV9JrFVp0IgRdNp5mShamb4HjPRTu+Wrm3XpQyBP/1Cc8jM16P7iBy
SWnGr18W8IgSWg8EWgdr80VXYFVFsL3xXY/KYIYMYl3cu3ShvZg4JeQx9WGoJBj8VlRccREqFW1x
//8EQtayT31rP7AaMYRroLyedPdKp2IU+NniDNMbqu7EpVfbIJNbw+15GDrM3t6rVN7xMxeH7x3s
N/k9iMeyaiqEegD4R8iRdU4GjdjpYZqE2esJIXYsU19teObt40JnNyT54Uor8c+o6mln81Oe/6kc
Emlm+FYqE0Y6yfVBQP2VbOQonuZldXf0BFTSUAXAzcmh3yc/yZbe5+dneDuklpgKHSW93+cEvo3B
SQrnisQjD/2qzvX3D/kO2DO36mZM4qSTAjHhKn80TXrypX/cuPKN/KhOyRcYeg/mr0xHZRM9Y8x9
rgLzbVK24RixkykAJ8v3/xT24aKqxaw2f6YL0lHAimg7koOVcdpMD8gjOz6fUPt0YEsPUHnsvpL7
Af2z+ejrsL3xSMkkJGjfeVeypHWUfUySbULWzUFc1PHxXvBqrziWRLsgdIi2qK1GfUTyGkhavxbJ
K+qKXRllAQEA/QSTUocvNNsSV0MAje1ucTvE6nbFYrit4L1UfNHb7JcH5ap/CjR0/B6I1iKyWT8j
zkJYjWXrjTtgbVHNS0tLjcLjEiuoGZ7lg8UUEQJ4CvLx2mkJVwkT8IUIls/fux4mv6MUpLqmHLsG
NfARmO0xqrThND3RBg+Yv04pp3YtuHU+NcVchHkmi7JrbScP9xWu24xgLp6nJxhFMn8ck+fRxU0B
Zp3kfvhsOpp3EjHV/y1DJRWwYEthkbA7DG4dZ9Lm1RKgl2bCxQHO67vB5s3xax7XA08apTyggmJz
fjXKz+i4evbo2FL+HpvN9xb1+LXX8zM8Od7FNUwH7a4fttLR6ZzGqlOL/yAyl0YWE6EIhIvJUbVK
WxjBlyKArrAUrSxSYS+om8TFpmRN6Rc8LV8UqDbhoYk/yhVqLEUjVUPfgs8NeMuNbWGdWTMfFVfj
EMP3qp9sEoYbFiKNdvLmu5jAWUYoEVXBMWqb+gtubDBzas4N+qr6ZeSQKL4fvuJ9iXx7vPJwLDoX
R85o+UToUcmyJI8wTr1ZJyk19CDSQsZk4NVyCrMEhv59MAizLtqiooQn0tAScSGL17ocYvGTRrr1
nScTBvg9OXl4kbjMIFWsGmGlHpABMk/VJUWCVKsJDT19uc+5T4WTEKqKmIyk5bk4Aj+wZFelxrOW
g9ZuZXom8OZqUTlrhPCKcMDBMtD4JPMbg9ZV3eAUpnVq3mMXFGu2R2P2eNNErvVHyoPjUgWLrCeX
rHs2AA8o8/K30Qc+lINJdd1N+pH3dgdX2Q4S6kohqBpzz5rF3K2IcIHq3IkL41x2Iw7mmDkKfRjE
kURN+XkVioCNs+k+4r1bMuaLTwwdoH1iZyVtT8pq6OgRS/B1fbx1UncQ8CaX95GAE6ZHyiqZOJX6
P2plNRO9dIcQqHDQREi84Pvzr2RZJ7x71SIF+pyplhzdorp1oFPIX8k58ISFBmEVnskzFP03Y6lO
kxT1kCXBbZOAjbDifSHDT/chm4WYu44YIfykuoG58d5C/Px/kfQWYh0tjhMPYwOP0nbY7YsmI0Jn
BtdSlNtbe3AUdtjiI6mxsYdrFZDPMwO0BnvGTdhu/q2HTmcYR9Mp/SIiw8+be08yCtp5gLglCF5d
0UdjAejNF+pU9k7L9ygxj29wXy6IBB9H5nWaZP4GyH9FfR6w8LbX0hF1polJ/MfwqORhRrqPR9pQ
3MtvZNuZA4em94KNQNBoMX2+7s+RgaQpVG54lm6SEfgJPxinsevQpfp8Wjb8HFuz8hqdgVTiEGX4
VK17g6QiEHuNP/LJTRokP6Y9vpBpTGEzHPHe4rCTmIMAgR2fK8/GthI8OX1ykv84YAVfyE12TCkU
Pgh4rejyx4allbO3i5Os3VflQmvwBNEwSE45PZFko5PvzK2PWeSfzVeEr921+2hbTG9b4n5BEPzq
5T28XmdTvF5rc2GcmXMMIbvGhVB+/dkyvPqlGoABxW0wMKrwvGfVT/cLO6g3RdZ3Ocq+d/JZb6z5
z963Jn/eg+YA7Fk9knYmMjsOq4gSgUqX/C9sDfJ1yGreVeO9LUeD+OKNZuNa3AaEYVn9JC6ECCxm
LBGVtna3eWT/gLet4ZMTZkDngxv68uuyABLCMSurI1S+c5dTLdZ+BpPjgAJdqclhIKQ4nPImzMra
tfUYmIBZhzvF+dFrYEqTATNfXrgM2jKTWVjDb+8xJ96EJZsV4YMjnfJA5lcC/7mbk8L/tzkdh9Ul
P6RnfWiMPZkQfNJpmONdIidltr0Hv9ZVqLVUpxrEyGOr5Tyo0M7NHZcXcX+dNc3RQCT8hp8mLsUq
oOUfiD7NXiuJCGNP8xeh1g/nSezMfcuOx3gzzn7U317E0VDec9+XoHL6NvxxP7mHmDFuwHWt+Wfw
3JJhv+1w9wazRncNAwwTeETFWXk8nxYuu7sULY0KdhjMdhZPNzGhInH+ZIcDOwEsnrZhmIaqdj5e
JTZIXaIApvhJDALeifAAPpljngKGhaCyoBZSJGCDxGOND541aq1yJnGenLkvlRTxdaJgFGDdH0XJ
8TchNKtSh7p6IgRzwodRz6PQWPtnRfPWioPF5Lxoqd5xa0VNmee+N8y8cC1uYylN3TD0mAU+Fo/i
I7tPV6yN7A610827mHti1C3o6e6+CXfelBk2e7koZUmnECCTgpZWLTjjOVAGM9DzMRpehzIGprAC
KdP7n9BY9iU5kYB+R/CGipkgFaxI3OiuEkgbhQJ4raUA/RR9+GljgYQkdmKlEQ3v3ttm/HpZjsmD
D9hP2+fBUWIk2X1EoZ3sPVwCtEK9A6HQDJ6/QBGQvGaqTZNFYaNYvrYllU8M+sk5UzwrTDuFhcKB
dxxTAUc6GTxOHqzMU0VlD3HqL3frnNhGJCRI+MMyZX7rH6NYOqfJTkOhHfOB8kv0DqM8M9Y8dE2x
ilGlH8tlqs+8eHdW/uLlUcT941uGZ62p/4HWmFSBTn+5EKpyGT15AX8DzFVJ7wqKs9yb9BvmHEmN
ilk5dWi6xStv9ZpmsYD/dsO9rfmAgbgbz3icp+oGzjtTf45qU+yIvFFOHkJ3XdYj+shSuXduiEp3
w+8Wob66cebSzRCvMgp79lNFyUL8p9SFlJjeiHpbxwnpawtjTwF+svRBAiZTcEl31OTeYdQnPUhk
L7UYz7NdxfLg1MjiYStRx/fitmmTn+ebIcmXfr+nEjardLjzPkY30ofO/Mv7FK8CWvzvsAkBE5hL
QnmiPNfYL+gFi+LIfhQU9qZzwyL8u0ZJbDLnl7bfvN/ax8gXtITJ5WEaQIu7bjaNvUway3LgBH68
wCjfnkaOjkvTrkT+enEkpTIhxNh/I7MK4rXJx1j+2lciV097xBrhFiyfL4OgEHgOHI+TXPj/do0v
1+oFyVI5KcSfWxsPKnc7VSojfTTMAOJyFRo3KvgIxyGTRpuM+SE+NaHFwhl3Gid2SFSAG+fyCjOd
H/Xd4NPZFOkQrjlnkPoEqr6fSOG17p79eRrav5h5fL3/S+/Htf0QsAg3JJphM5n9MFpR0sM2X26M
EynaTkQ40XmZUtoWPBAotEzdqt56uC9XqcikhUdMplSUT5uXBOXFH6bpO3JP9BBS4rriBSkC6SHO
2FFeYNlkPpi1/tkuSgFYI2g8dvyQsTCmsCjZQi29oHlHOGMyOcHCjMtoS1mHDKb/cXKtNUZUod8C
chqONS9Cgh0SEbtHMx/lM12SW7w6jge6A8P0tZecnLz8nbGdXjLl3hUqoVCmAZnS7k7QiEXtSeLk
vL5yoR5gzlFw6f2Dt7wP5/5/PyhPYHRklgrGDuRegp7OnJpnxEkkCao93QgMIKbGQHf0jJ9ImaGr
RnDYJa6lN4NH2FCaOrA6PkG0ZSvVe7zmPvs65kqyYzN7LcaromIZZDBdo8TliWv3sq0FhAHOPWLs
ceD8uRY5CML+8fqusH9bNJRcqcdErKLGYmksuW9QATaodT27vdqXbukcN2lgzyGDCFz5GhkQnxPW
D85dRTuyJ99fDhRGmwCM1m8pPqD2bqWh2C53V8aZZNrxHsBC2O6ZYUDabx/z8d+0WjMQGI+joMyr
oQ3FTXcGVeKjzxVXMRh/YLAYtTHafTgviFlGOmmXXPN+jsbTnYOAVnEx5gqWzeWwYyzfwGza3jOO
ftlz4kzwl9r/qI3fnAytSKAvguiQnuHCQ+hbOSNf/QZHTwWEVOA+DseuS1mH8gkMLDrAK/iLO9IB
BtyH2Yn/ETkEbNQxlbLU6i4EfSvfJhvT2ttqMNBJSFFuqNyH+ZoLtjy4LUIiqUXfQNvxruoUIIuK
Mv17lAB/NRb8/8065QtESuLPVGdLoVQMtkFXWnHkMcRS4gIafcVjAhc9PavSpPSW1RYHO+zQ7lfE
x26vvFGgoBkxsX5J/zIhyRjxzuyvukC/nKGqkM8HDLFFjBqdim868RXzQu1WgIMReB3JpSIRhXKw
t267XEvfo08s0h+gYay3yz95uHbdT5YdoUz2m2FYDnHE4lom6cMM8oZmxhVQUVWXNRDmwsHyCRlw
QvtJ5fi6xKQjfJ63QTW2XORpDLvWBjs+Ydnnln9LZIhlAGufnHv8v+mHMYdjKMKxUdwfE2/uxsdy
AEFkG3kzBODD0jzAZZuSsc/mac5v64pOyBiOBQlz1YpFYu4tbC5S3vX4rkTgB6Pho9ppFFUuAMCU
ITXeAgbfrpfgxwTpIRPDDXlDGIAb9XwrwM+V5gQwMBafZYwMIIl69jiFVQS6xMTSSNpGQhRhQKj8
s/OJM1iF9kI+ZGDhJJxVhKZrfmKt2y3R8MV65p4sj1D5NTPAn3Or1gNbm28hQqaiZkB454a+F54i
7wcisx55UWOJ9bZj+uWEYC/NYVEKHBnExsCKUjexqHlzFYGqXpXvz6uHC4+gH3bGAa0E2KPJIbtf
p+v9xF4y/s/bHPI9D4WLeCpmXpOk0kKfhUlUP/aejKZ5r0H4Xj9IrJQcxonf2XQaUX6Wn9YjHjEE
gZOcA3WWvNc/oY7bJlgJGTj5XUCgh+FgpsRujFriFGwjYgDsOZLMWpZFL5vDyLrRnaHwkBJkayk/
ivrnUJl0nzWSDgp0oMiUNPa1deFdURQgnh/tjSvRkhx2vFmTI02aRixU7bnkQsmbUwY5n5qMpIai
OVeXY/fcgp+wCpHH8rswo8+6QKlQGZVTbA5+1VAMQM/ntHkm9vjhNN3CqC9j4aFq9kkcmqwuM+/W
KoNxViyN5GUT8B1Z5pH9G7ODfF+dSLlEjNqidyAdrbAxVY58tze9zaXW1LkPWIQp1uZRolGJdndK
JqObeou6z/Yd9FiZP3ZWMkVLE+zqwn/KNJixi80pneoeD682Nf5/JJ6gqQdAEW56Zvj3djCwOuhz
hBqDdZ3eIRbiR5EuDYBDyNzNALt/t3HJeOBtRWJFkrXx7LGcpLvax8z4fndHCYWy+VxH9nSiFjPx
+HEplt8gwLcS64OOOUft/qDOihsNeR8Ey1OkdHBiMCLuPjbBSbvSCHl2qrNFjMzW4RNQdBK6+es8
j8a1H2yO9uMFlWvVPQRPIOf/AaAPijp1A17ukjlEho4QLDelXNkmMQHxeoDmH+83T8U0CnYlLbQ/
xJDiJMKFMnh1N6wB6ShuDCZoNSYDmB2j8oWFSXKheb5oi3YT3Mj1aVof7LqOx9LKtqjMLyjOXWfq
LKA3QIye0/GfuaIYHoA7WVkQ2acV8fy7vZqho9IGnMd1Uc3Ah7Ry1uqM3ecld8IfifaDfsS/e+M7
qhmZXnGu1e3C7CDnHWSeFWIT2n49IgRK242DG35k/rc0+Z4jx5NYTDHRfX4a4qWdxIFNDhYQXCtI
2Ra35Zgx6N2xgJe/9g3ArUdvDNlktvu3yDebaUrVmL6j0ojYexQ4zj9kDqVDSu2zXpKcLDLon0AJ
Koecw5xPScs/u3UmY59rIG3oX+CPAdjT8seY6AfsDrXtErpP6FQbVTh1RalSHJ71/7eXsTGfdOEk
7ssJs+CYSYe06twX99xFRFZzdiyBv7FLX4ivyW215zVJnwtgbqBxXcr/R1/zanbdAkU9ShN5Kfp2
Dq5Kk1Uo5H+eOiafltXucGmmLxSRM3b12JKUhQNjegx1DW/sIs88Qoq5+sSKhew1qWFymTd0S8FS
km7VcqyoIuYD0QJfY2b5RGl6gBNYJT8WBYc4gxlpe85RwniPi8Q8EqKuVJh2d4nIW+UOoKstc1PC
JYatJv36xeAOIizre141m7fbv6u/ZW38vMWlLxxH7rpXxtl4ZpaGxwnRnGAF71BE5zAb4B0IVth7
l7W/ssowS7txC+rQ1ik9pCEBXbGw0hyB2Hq5d5TBas301mg0hPxATWPNwLQumQe75O7izPbGRu5g
vgqR/HcagkrtYzYlxxlUxuRagq9oZOqTu8PZDsKodHFR/gghEwigOUpAtLS9umwg5i65MM6bey7F
SH5KQBLB6J8xFUsb0O70sQ/E0Ee26hRSzRlLzkGrc2kJ5oicZpvxrgo3LLTMY00MIS061lA5Ytnk
KmmsBrrbv1KtpTbzsLh8Gd4C1rMFj3MaY2FqV29Au8cuUhkVYao6KFmGZj4RKDDCfGTYV5db/nSV
ISmOWC5PUGXivjktTYb7/a0OXyu2N/4Y+VkUK5hBMIV3nzfRJBjDW46K/ykuXVWYIKwpkAhhk62Z
naAHqDSmN4shge2iLpP+waLFBVES5HdnNVVtPDY4AOoDtwB0nlMmkMlT84GrsLrTvrrr7Lve8cB8
3ISzK2xsh5C97dBXl9ifyDyxTHyVLxKgatQp5xg7D/S/RxP8k+QZDlV53qhquOWVcqWitXQOgz6i
3lwaevbtOchfqcrzztJw3WkhFWXskNEcxNVkmOZC8yDVjl9o1i2CGgVvWrwZmoo2olH8fQMwqG7I
skE8UJqIG8EhZHWDFIFCFM3nHJbAU12eAKMFg+TNSiwmzupI8uTdsz1+sQaC6zTFXkVkMwntKcTq
AAT+0lCrU6UhqTizRQsK8brYJQKt/b20Rc8XYcIv5zODjYViLuHtwzTl2VmKBzKPDhkGrO3NO4Fp
JwPGh+QRTQwe2UN53AXbXt54rGLgd3DM60LtbI6xoJze0yBkPbhtvwU1BFSQcDQlNUXUWSEwP9NX
ShPGtIEeaX5UCE2rmCvvcP+ABdahI/WuELmWl1fu1KPFWwKYxwNcFBZ/2xJUcuTuRqUAquciaFVv
gqjDPWvGkeCeeOlngX5ZaYuPcXhjLaorou5b/4waDO50gQn45AZhCWKw+qQMYgSFO3eMdN5PU/0H
oZ+xCpz/bjdB2TNLRFhqF05TjSLD/goKFxBl78XiSletGCRlyZU8rkLm8b4o2UTiP/4R1H41Jppd
24kvtTSlCNgmuGAETyiLL2+cSKLwtdm7aEAKgmcs8kM+kg3o4Za55iv9kBqMUgfB4dCxuCcxTj8g
DkXo7RjiP3byQOky/YYWfKoRqDc6egi6DYt2QgpUzmuI9Z5yQ8SW4ayGaj2P9UzLp1Q3CdMi828C
AxJ3jPe9OpMHVznzr8Z67f8wN5FY1A41DpgOdSARqxgxvMqUzbge9cyTp70K14jt1ETtgNEaC+MM
nCi7iWOEaL/TyAnm4SRW3UhZdqPZA99+yoFBuydObTMIzLPn2vN6KlaqmyUlajHce5Sn7Q9RYOyE
2daBJKo0yPU0HQZc4dy+gvHGh6RJ+zHn3HGKN+pF8ZWBvgJ0NUW7eYS9RkB8tjlNl3/61M/1lxYL
7IcznnhgI3VjwWsKWIRIkpBFA3EGEH+QWaqI/i1RF5USEiVU6MAwSDEm50JForHIMqN5Un7arqsi
/230EbeDm1p3c7h9rK67skf0+5D0qgjYpbFF5t6O6vSGf60WZOkU/ZN7kyadepmbkK3nPwxvBPe+
6DaehYoKtqRDWutRIIFylqXrvo+xInngS3Ols+yal7+Qs4C++6g6KM+mKIqp04j7XJnkbX0gCvFN
c2oXFpOtQIzdCbv9xyW+k0+44JBam47E4dXVd4meXyBUoL2AvFn0Qlzj4L6JlCqVESjiV+jixOaT
LtvYWf7K4wJ+RT59B7exzP3K1bClbE+SNdqueADE6ImxfOMbm86faiE6G7sHcl7YzM8xSsFMp8jx
P8m2JLx+v7gn35hOC3Hux49/Cx9/cSVfflefWANhPtMKiBucEZZLcmlUUOZ0mQId+010040iJD3U
ol0M+E8KWTwKu5Bf8C9uh9Jalq9fXfBy5BPCS+qdgGJibx1ZuFrQ5Cf95bWl9bUqyn0JKTpmigHa
gs4o8gIA0wUlxp3gbagBz88u8nX1wL31+6B33PAvAbXYoT/p0P1qgUyNbxav52DfJ0jYOKYlGsr3
i6/z02UYmIfoO96Kl7NtwRkrDxHka1r+iCnmJlLVFrQ0i04Jn7yh7Mz/FQB88XZ1ykMkgNxgXU68
aaMmoZrqsx+iqd2V420PZXYkAvH/IVDYzaagmuVxV3qgFhkweCYq3k/6bRhXXuXQtBZa/+L3bmhd
C6QU7spOkBxWoSP6SUFhCagVGOxvheMgn3tCn0sXoXhCG8puxeBLvZvyYjqsqHH80cQnhecMGfEm
XvBfYzPchAa7ua2OE+Fa6ujiHs9XOkc+YVdo/zG9AL3wwq09ecAci0vj/5aF9D4qPI9Ed3MTqvcQ
0eY5XPHszkLrwtjkDcHQB3Tq+IfsuWUC6g58JtsqXLzTeb3oYDwTenBk+mXXzid7UKDLNu4QKYM4
JSeCSrNg3rV4UeFd231MNUVyF5T44ooEWq+PaeVOQFv/N0vZjyIblUjsy1/cT1rZJaOh376uXHf2
tY2UdXYac9WjDhbSi/zsrWNY1+jNaTanx68g5mIX2wiDVted3VIdQ1/o5Svstd7eWxyS3qqcYNbm
jfRW8E3bPKZztuvm/ZuP/73CPxaXet7R2ISgcB8Lxwoj/ULAg5qB2AUKcympgcJDJvoRfhi+XaZJ
vC1HlGWmTfHc+8s7nc1cv0pSPkTVc5HKtIdPkUu62rVb2N96zbOanOIaOugfIStUJZ++lV2pJbQ1
8KX03VjybtbThCyq1TCdwmmxL7yoFDWeiTVpgolMvr9FbM9/O/0QogwQ695NAsl4KVsEjhmyhjS2
6TmV5tdYBtg9BFDCY2USIjNE6M03IAzqqGaGeK9c4FAg98fVLvt9+NRiXsR98SNmhOnVJF0OdHYK
D6e8u91AXwpuGUtnEJzkfzIuSXzJ3WlS8VBoBfAXiqBIZwY22w2V/N357HyE5SI217MeJryZ0UEp
+eDwmROmUg169ZqmElps8dQ24MjjiJ+CepuhDfIpJNTvoagtwi84ArAwbhf1XoZ2KATabe3OvX/1
Z/fdOh6Z5eJ7e40EhCYiJ30Rtmk1WGS0Ee1v6RaAukknvjulF5VeBvu06QfavSemb45DyeUZHGXv
X4wwYSoh5kUtE5TrUd0R4c/D6Ip74qociWZX9TpuKmfoNjiC/5cokcQ5jVEqzCHTKE/aADIuQ47L
Bvw55tXLQeNmSPkF5fwcb/nu6c3YAfHfqO8Zei2jrIGOe6f0LL+8j0kmOOa6w87ys0C86Y7W2NWF
PsBo/kcjnIsumzfsXT1cMZ6lH2fFEa3uYxtDPsp92kCVJ+v8u/28Ocdu5Ro0GlS8eHnJszrlhcAR
i70UGAUt4/v4PerPGwEMMiJziu47LmgYUopOO1XW0tF3lsvjcFaJDoOR33yz1PIxg/+Fl7h/P7Yt
SjYHpkyFCtZ4EVa/tZ40ETwyDVWEcBbXLUeDL6L6YYEveg1YfxK2zPMCO5//1haRA28OZskONSyi
GBnOaUQ531UA+g0EgIognbE6DBHBp9kIwOrr2KLnmctKON3anZPR7GhYgDz83KG94hyM3Yo/9WbZ
fLSEBk3xC9Kwg91Z6Q28janwHZtLspm5XdCOaPUPlcKnm6wy6JCfvukXiPqXC4v/2k5BZIb3Anek
4aGg17ipESHcP3r2AlR4n1xUHI2IfC+nm5cXAOBnfxXq68Q0gzMRJAsyXNQ86+k6MAC1+YHFeJTD
1KkLiLUvfe+Cbes+xQbout+nfpmb9UK3G02uKgaAKmUH1PpXz6gMRlyfp5t4qd3bWPjqgMN6Gz3n
Q1JeebrZUHqgSO2kA6KSlw9nkiOlqy6Eo69YTFaliIY+FPCZmc8Ow2vn6vuFy7Z9V7qA2r9XakHX
LHmbTEuB5BaWDoMww+XruYsUzNg6Bs9fz8S0IcBEuxmkbJl/us5/O7sjLdeqxgzyHl9bedAVYYUR
LtMG0FsoVBTTU9cOz4mJQcsYxMW+RgKRrZxSPvwdOUD4YFwel0kagYfl47OdTkulW0Uqxgw4UJZe
jASc/3/jv24x5O/8+U7sBBiHEl9xvj25VoCSXWXjCgFkO41daaaCq2YVvjmWYlVWBXbCnPZOMhWB
DnpJr/qhzUk8R5EDbQREH6i+3u2NIYwmVCD1scJ2U5qgkaFKZAai/GI4Ohzq/4qsd3jo1b8f4DVo
viO9wOo2cgz4fa/G3ndORKJ3YYskhCCKfnMylb8Pj23s3NXKp5O85XknhGgeT/bRe70oR5aWCe5q
z5umwauBTt6i2pvuFRXuDiwih4gKBP2kngjUL63uFraZyz2l3zUpzK7xvNFV6LtAM6ZA0nZhsiYd
IYxkKHMKRrjSiRHF0gBcE0qXn5N5aZrNQHEV7Q10j2aywVUsqr+JOufV8dT2gNIyQg/WrSvF3ptH
8QIVFfGqKO28lafTMj+C88sXpPoDQZxU2v+6feI3qJzEg4r96pWInYEPybkOYHtxpicyC6k/kjvR
DIurix4bkpQ4XMz28rcZUmBvbEjWFaW6cNm0HEIJpqV2VWcXJWphUppOSDrbyTgSuIH8X3AoYSgB
2MIVhHkrzi/uABfQRcu+DP6oHBZcau7h0MoGvMBcUlYdWeYD5GyELdEaoMXMVu1mZNgoTMKj9NY/
lXwYizaP1h5GruY4eM5pRgoJXMrkc8QVScsQTLL9mEnZD+FPEvd0yh5sNyH3+WUcUbr+0qbS5p+r
CrtZ61uruKkgJgmKnZA8xmSrmKnpLZPvhgmP7O39xWckMx9u9ik2XJDtCPC7eupFSJ/+agJSg2Fe
2NgPgipBVW/n0GOxuvxpOnXKWIApkx6gzuZOvN/62MNTTm/k9Ss13A3KLtOu5Khw2KhrsGmQlmQe
gy0qcpOXu4S/quN7pazXM7f6RrrtHRuWAjghwN6Yw8ieBw9TBMGkryg6V5Sp2szMUBfb371ZGvc0
Sb789xNvcAEUAXN6NyAL1e3S5W+z/W0/6Ll4iMBY8kLrzpH7k+ClG/yl35NohraqJgXB+NFXg9rE
oxXnkZctaHQiIMWvlMnDJPM5lg8P0CLfo0j4jPNJ96kTm9ya5EJHX0fss/0KJW4h1kNaickS51iB
11z4YPDwEmWuLFbualjsE/W8E8MEhWihNWQ6R4fcj2WKccUKy6BU4dLqn+1TMc3q8ygyVTCtLoOT
9o4Pq9dL4IOWNiMwjtNafp+es6smSN5VGTwiZQ2reP3ShQxB415IHGFjKL7x5lVoAnvX8kIvK1OH
ms3FiXzX5hEb77o1VHjgeDNOcTxZQth0IOsOaMeJeVJS6IUwM8Isf6zMQfAhRMlG5cQ0ELtl5Jfj
XsmlA/4Tx2/yEUn6PMLhO4eRT6z/4K8RrDa7BEFJnVKW2z6Drd5wmEofxrqOfg/zJu5+2yrBOtzL
mErCVs6F1EGGe5rJPYdegaTWVjhvgDCDX6mAqtck36oUw8IHs436YVM1AI3YrUDsEiAT3Cxh/t0Q
0t5dqIx00lH9gkv51UubqES5Muz2mrXyJr61PmljdqFWhR5/OD0iQal061XFb9O5mvymtjlaAQsC
fnYRgSPgp43mYKR6sYhdXeJAho6pO7emBgDzAxLjAiK9v4L0pUZ/7NedY4dWDL/ENvwAZxQBTILz
KTGSpcAV5XbG7r8fplp6RcrEexm5h7VSzvx+260+MXafdBwFLyVdvuXEbIW5hBk89E6sOaY3nSJi
FOCFOGQ2EoOZN/mblTE6OtHBnT1B47i2ZSifJ558rhmBvtdEQr4xmA8EuuLebzzOPN1b/UaOMDzY
wYw5ca93ntgswdYLx3CWY0ZZ1TtMszoiW/twbny8wELiQrK9Hj5C2HSIvT6iqQ8JQibn4XOni79z
FF1Oi1Kxd4jXGeznXpRwFC+uwJ4eBWwqxcOatBbXW/xx/ZQyO2il4RzEx7h/Y8Ms5ZRWTNW8bEoy
NdLz8NTnlm3SDwxf65NXLqSv+z+DHKe+0eFtpCrNHUWTp0b2oIRgIL2FAFKuILxdl9NW4raxDboa
nNj0qJdmz0at50DG1MenWinlcO3B+kA7GnvwjZ8qi3k+AcdJP1l/7g0tlJSz7KGGgOkr4mJK6MBs
ivsu+0OLxfaKfuY9tZNRi4ycC5UTpCGZ3ofxWc5dVeVbOmAXGfMCc2muNX4EZVj995DCF0kgIHys
rIccAKaB6DRLFPCl90k7DrHdHJcK5TX+X9AzlPChit5udB6Dl5ZDAd/+3vAUBFoaXkynYkw9eulM
8YLv82FOR633rWbtFAs+9T7w6RDE2TWCRa7+t2iawYtjOhTjdbZMgfK3htFTJBMeE8lpq+NAp1Xv
ktgDf7Wdas2JVCiUl0y5czn+vJJUqpVRvFl8EqpeTA+o2baoZhAD1wh7K3YOS34k+6LhPL7nZrD9
jea29mPUHymEehhBbaMDMelQCGrLl2xMZatdJ1nkdxBeYtRsZ6Bb0861Uka3XFj7Unv90574T6A5
h9CYtx82GcvsPXOvVOYbSc9AWsvzU5/SIem8SQteXGgb67XyC5UWPFIcFSfHV/dnGGuhd8KOAYr6
PIIbryPPyrXltIHW4ePsHOrHgSLx+aEFAyhrAOtS9R2XCn2Ifb3SHpzjyhcJfexRFlzRMqaHhCg5
U96gazkY+dkNe2Il8O90yjBvT4BXRi2+4Uv3/vjFaE6C1MWdnASW7m4wy7b5n+vuN/8b0wCzejuR
p8j0v/uzff8zGpNXELqoNKRz7tCxzGlhj/ZhvROdpU0jtFudoNPzis4tAeqL8WpZxe2TtQgnwism
/bZ2vEelugaPUwdFpElkGMOlm0zONrMKYLLmD853jU+O1NOjFt530NbGKufFL0i1n1nwjb2KVIr1
oR6JUZsS2FWLn59531YUZSqIWH3TSUROP9NOLWAmcD6d/ohdcofT4kXykOoXq6CrEEEBlqZxd9Tn
ifXDIlrGLZFPq+SImlil+Prl/I0bEbHZzDXDOB2DMuWTsGZnBnwmK/mxIImAJRcYqe32OrGtRJqu
FBkMe5crc5Td46GvcSXifdQj3OdDyVw5lcKEOUNtrnCQz8jOyZJnajCiAiUcVkQu3iHjKiTd+lPL
Uxrts6kmasO8y8CWrwTSZ05IP6no4I+yrJ8viMurbzj9OKo6jI6+HVuSItcAQXGXfOZStHOb8Da8
cotuouyLonJ3gbaGQ26czzZ7Np729X3QFhbeth9bQw3GRXsZFjzayMpZS4G1IsbNBvWtSMC4LBkE
GFtC9pG1i3DhTAXKFXmYhiB6bc/reYv+ZBQiX3hwC+/mnCDqStjwg2razzKrXAlss0xdJsdDhHXc
CiqUF4k/n8cHXN8r1QaMx29Suu/SzSZrNaoSPasJT6R5bRa9/AiazqNWpohaPJFOkhfIDa9I6jD/
kgNt2rsEheV98qw7vcFuZpnnDxWH9U742CVPjUa2PJ5CDswkb67oId2nEPmc2gorZ1lvOZ9FQ62X
yuV/hC4+Lbt/rTuWOBst9KXi1/f1qJOdCA7+IfrWK/pl9yHxlpOk3HSIUwZVd0sz1QdUswjJXqIF
i8keLNyD2rHOwUlzfvdyAYXFTrJn0XS7V4CmCxzDOf0d0wt0efWq5FYcuPbWJt1XlnBYTh713I9M
Z/p4tDBgAFqOYyEfO961poBWLxkNdvDR1iteuy+pPpisfPgPw3asGgBawVfzmXzRhBYOY/Qh4V1C
J62xq+IySu5JExHdmGvN2wM90PrJ9cSfzZMMUtVCEuS7DTLrCa9NX67ZpDrskskKsTvOwPAY0Z58
0awysA/yJLAnfcAT0bf/gh20imv6ivnL4MH6iRIEdxLLEKlN3oygzANiQCOlJAmyETzeRtKyjP0F
PAYoUAzFmGUoEyWWkVPqYYCaq4E0VqvgnriCWtZd8T6CQoXoJcdJAPIxWTv83VUvVSptawXPvYB3
E7ttzMy9pRGZKzaJK9WC36OvnVxwf9o5LeJ9RwpOVYbdcjP7t49k8vig8gxvgsEsS29v4QXnRlIX
DXuhBNGfCXBthw9ejVWzJsKaZKPVIM2BotOEZnc5m4T+J+u4Fa866uyUHOHBPgBx1iIcIftPotDV
KKgQSF4ESfYZyWVUY6aF8QnoIk76qr13G8FrishQTjE7eVzjdrpGcyt0ZDjz+93sAfBw4DMptTY1
02MKaXGZKqjEz9715YadZap66+PWmZ0ecrCpcRTJaVP0YuOXh4BcYX9uRkLZMm/CUQKulm6GT1KO
uwOWcmtr+n9a0q/4zCUmJTxRMG04yoiVC/ZeaWFN6IVl8ThnN2oQDZ6VtsorIf5un1IESgWPlKsT
6VeTs2GnoX+vstuID9/5ODMXRl5UUR00zpIJeZXShjpaDkxABl6OYvYXoHdjcMHp/btOVbWBGpex
pAxb3irmHtyordD2/MfGii43sN9HZLT1yXrfDR/bRUq+1nfsWHLV22C3ourTzHYWqJBC0CE9174y
uFynSY37oDUe0G+GrsaMwToycTGYXwO0imdqiSy+yXn5wOQSS6P+VsG3bxlnta8ltktLf2uU13OH
HYo8omzXm+I3UZcdBhzl1BD3g/PJrgw/wx4XD1vNnBKoSgZKnpI8hGDP6nZzD3+0LSTkfqmmy5gC
T7HMCUZAPCnAhm93UOHDSvneVMsUMTwOgDiwB/IFnAL1co2ybVEpoagu07fj2PGWwSNzZOqkWq4U
iDnnVTeuPYL1gVSJO6QWThSTW1/v30S23leh0mvs0KhynXLlQoqXB9JBgkNLz+gb/ns/mvpJMOzB
OWx/hvVoRV6Maog2BCxdVhacJvwLFxLV4LmBnftbmY0Ng/GED+bN/1Wy39K2uNkAou/QldsuPsBh
qwvf68rAFkmsvjo5w38Kud2VSKM2PcCAZq4Xn9A2svmwVGxVa1EQv+Zy7cfNojIjORvUvdGbGKo3
GfZIfLezbeFiLuY3vzvePYtQvy1gIw+IuGdqA0fxau9dEouAGpc0hjmbVAKCGeOsnEZeqveSTf1d
sy5kMFu317oehZ72tUF6Ta5ZWiETMoPXZiOp2MPf3Mdp17dnvCjnpCwT6jVU8EMnYmuEH1Xr4qAR
BuS1G/cGMmlM58JopdCwGgAT82Ou6SsejAYO1SOAmpZVm8+1l/02tL5lGDOveloUuoSMhJmjhqa9
KbVnMZxr9/fzCkEh5VjdAQrgpnAAPWtdlILlpYDTWKP3aTM662SN1H+mL+v42tNEUTIAyLt1dGou
Ih9DXrrbYkg0SElqQ2IpQDe/8OSXPsxYvZMQpk1BQ9DQCs4mW5HsSPugZiIMEAhIRNFjwFoyz76L
BiL7ng5WOQamSq5lrlhJ4YI8TpUfOsRTQJxNRH4BfDeezm/FZnizcgoLiHS4VseaEGD/RWEsCVFu
rIPYy1XenQTHqzAHXXt6SDApDeNvm1SoUw8+kXEvIha0JJ+vgkTbFkZ/z6WJAN4axV7V5R4VzOil
j0CNyuEOy6Z9Z2lziG0UxLN887TNVzw/UYO15iUegOVkosd2pzLvI3+AgFx+rePgwSawqvmucRIJ
tP/KM7j40cQDCgdm1PrcNcIrQ0hgEE1o8xYOvHYOR1aeY38wG1RuJblwQv74RVcveZt0HVF2Ei2n
o9sFCBJWbYkfzL3MNnGaJWi4/2Yt+DJ3aU5FNNsNzoHWi+tIo/8hoEDjmlDKboEqJH56/lUbaxih
N+iGTk1xnbNeHaDVPdo8jMyOk1wiojgRpvgO0H6uzHYdGqHj3Cp9tTbjfAS+/yw9YVuic3QDojue
bEIgiRML5yKOqkXv21imwkzm8oEe7rJBh2/zDMdqy0GwXviANGpDE2dUB0xWqThXVvpS32agkz+8
pU1pJ+h97q7eAcHpWCFh+MhD+ft29FtFpnpLT01GwibdT4RAAlyWUkQQXuQu2eYvohhFRxwV3An7
5roUbsdm78U404B1dkDfB14CCzUuqgeaYkYEZ0KbUAEjJCzLm93gP1BiSebsgKLcCHbXxTuMoSSL
0Zba+CAg3Ck+45E3bHmRfN6SMaFjSkkGPRhb7z/VfwSOaJW7LUVJvRLi/2Nt3iEPXmVAXL/aqU6M
rfal3sxcV0cHYOK4WorrsbDyoaNN5m1A+W9zWrb4ojel+cvzpIAqnJTuzuSStkQwSfXhBcmzbAR0
OoGJBcx/UOnzFd5TZnV7fxWv+TexfMICTJsTJbFbXGpzea/rObs3Dcn+/WwvjMJThPUAxuj3MysP
tdQPmmcBUySDoos21/tSnBKKSwkPu+3Zp7UzqAvxyiWke9h6/Y/en9tSZe8cwNGieBdjG1rLV5Hv
+Iwf0RHVlXOxADgHAsfl/eSyYTB9nQ0iWmKxYzOJruNpOPoXvpXubeAxYoKO8Diwx5f7tA+UaFLZ
blfhsxtV3DkgzGOLgww7bNzk/G2rQHNHQp1O/AXFkdISmRvOkNQLI19qwvymV42rI0NKbGTwVUym
qwEO9aYiMD17VtTzAAiBQSDO4bqanaLQ7mGHDP71BwbqzNVLajEpy2xMPxqr69jCxnMzKqk1d/uP
KCvwhAXgiBqDzk+kIS9ziiiO8e9om2mHhqdjgSMZI1YLEY/JABgzT4TIG0Xbr3UYsr6cThgARuNJ
/3UiEbBNb0iAmTOD/DMVg2t1MwWQoTCx2xBXie62LinvMEnEyVU5WYBeIqyuRR/ZoaJP9vgzvv6x
2mEJ2PKK2HNTifsObujlHiA/rMoHkBn4LRzpF6M6Aq4MLFleWmoW2MHCLd+BG2w9oHuPK7Smhyvx
CuKA10QzlamGcCYfeOLtR3yRM07cnAYwyNZJ+F1eAfSut8slHHUkWinbasfkCMK/mffqKURJqKOI
PXsRgeYigcSaDa4Ad868bNbHOQbVRdFEusOv+Arc/8tegQmnSPWDZORoDRCcz8yjekRREVfQmFjq
C7GHj/+kWLIOYdlqGm8BGhF0iu4ERkIcXcjUyotgyANadJiEUTYxU8GLH8dlRnBmR3/mVJJJ8RsM
/cEZgZMqtFyxTs4IPGC9xU7bDzNPvkPCUAnMxq85tKpO1URTVhTd1D+I/LR+8UjpdMI1TGvoUy7s
DV3tfushcdf0qdRmEhAV8enCN/H5Lx2rZsBkGsGkZlqmr37IiburbjFL+zkW/bVyoMNclvATfJWA
Pnv+sE6rghvdXH2JQzlNhPNFC7ETwKVWnpIU1fa0uS0bSruVK54bLxb4FXdXqg2PzPSSBsemGar0
kE5aJjadlTyia3VcZwAIc7idlXEApQtroFaMK+jeAh0M9bz1RYrp355IdTxDPax6rGzAskrIUcBj
8Nciifuc+jC+PMC75b1qQxV/qpSMzyKdJE6pnDbFA6XOx7P6rLlcN7W3fynm4f4IwDbIkbNAeGBr
uZ94fTRyHxPwLNhdZ5At38ftNnAabTLp/JtnYmEgJv3nIUxTFtg2UVur97kYp8VaSSQ0sYh4Xg5h
pxxPndQg4Y0AeMW5d7VHGcN6uWGISQTF1gKWiv3KjT1mZcavqM1/wcWbiDi+BYRchO9tw5Yb8JL8
aTBuEfORuD56EYBf0iesNkJiPP9UqeCaw63NobAUWX0qeMSxrtqIpZ42jlicNRXpwm0DlJOo5W4q
GUBDCO9A5cUal2PMm5DjA1k/4/Kuoqmc1G+dgwv/BS/ZghjzXOSXeLnoZCxoZjAxT2GEf7b+ze/j
SyKkMas5UFagMEj57hzB+VDufGR6CoLUaScebpMbgILZ4UFR48KqeDxG5xwViwEPoYlRffmnK/a2
VT7WN+he240giCddqxYOsnnnYp7gTkZQfIbVKDAj23A7Z+MgXEREc3DZc2CMkhFZuA4rqRGgQCzS
+2OYhSIiCae3A9j/4YRLAKc1y0PmQxcvur2KRLwbbCYOd6bVAPZmUAgmxrSkgWjBJ41wkM70Qqei
wGtaLhg2ATybMwVqtwGKYp9WYp7nTxK4eR9zByGurD0tibvYEuGyGqCszfCr0IMVegMx0Ri/hHtB
eryYKapXM/I5NDUt85tw8Gm335HqiqA03msRy7NQD2hXH0jj8BJIXST9NBEAdXi+Bzn9YRNTX5w1
dmcBYKrSGOVtcKo5xZf5BMegONROFcBErlLgKj6G9dokekXL3wdfTHindCYxU+xbN/rXh/YLLo94
LodjdwHi9L5UeLl/ZNQUAOMZ0EBjc0zy+8/1SF3gLiqxl+qlTBFwBbCdsJO11fCq20de+jo7Ck56
j/lee+0LecWFkeno23xjUWdkFGOG+GzLC7mtIhokpIq5o6q0YooouBlyIH7IrvVi80gWkN3HU+PD
hRpOOcNxPOjAwWCG54D0SufsQJR/ix9YBdebc5Ji1Fih1/yYgLxR8oof4v8SBOU/ZHP9QaMH1uef
dNlLql8JYmxYoYLiouwPU5IKJ8esvtAdmpbIRXx1ZO6FYGjg3vvRUes5RP6Ax7yuFuNxnuToyscG
uYC/8xEDUBSIttJkkchNmW6P+G6CMbVlQp10rEUwHymAgzk85gfcfkBk3Cd0Vb2SeIRNLHdBxX2s
RvwlokT4rjjMwJEtopJFihu0wxsInwaCFnPkUInHLUuicsPDopKaYh7KzzLE4ZtRXRoh1eSRTajc
tCK0Z4ZX3E8YSsqrCSriYpI8CREUpMdwyNjOcCmvbElGRp74Gc4rrRhIG9PIB8yGezeIhkzClb8h
5m32i2BxBCp7EkIkAtP9Zt9Rr2z05ubfhnzBi0fHZN6scs/DcT/rzKEBZuzgBIfwlIp819/CrK6z
W/zRLBLuhqB7hEvfg1Z4AMn1Lx0YsKVuaKNt9dProhNU6Ph5USFdegEhUDK/Q2gDODVH3Jb6vNSh
UKL05iRxeDT9gcWB3E5SmAmddUmeJUdn1fdI6uFMjp968y3rXLJUgRlF95dwZIWvp5iFciF/2pA2
9WccpZoS5icCFzuk0ElRcj7jxt3p3e0deddJo5TnDwRoU2U6YyZIKx2ITcq4eP39bCld8ZqT3kuq
TglI32GLf8UVEeBrlJChcrGX8Qv33+tmwx2v/T4B9XAm9gfji5pLUllP0WjgXwtaDQB329b4ZM+P
KtGP1PK+hvq6gXVWlVKv6aQoTidDsPthyEU9nwDXl0IgHuPvJbON+1nimtYGv0kkYtEn1EA/CtAj
SW/m+DhSAPoR4lt3Jq3oxRDlXutwH2Tm82Tq5jHoWmnVFEriyQlbvOP8MrAjwtOWnU1gq5Qk+PIE
HKpLrZouqxrtL1MXsm+BRGNp4idIv/IwUsc/V7LuwPZ6cdsNGa688GlAzUQBeMK3+DVxSUWy4aTr
zh4WffRmrgN3ri+SsV/aoNoY6UCqW6KDUbtD1Rsn3B7WQyEaAXFDpwPpm4OcP/AjsOY0FLTy2Bn8
9cWHgD6EByjX3/sweSdlvPNzS8YBSgz4ZVDHblaj6byupUN0IiGOlL/rTQGMwShV/LFNbS0XKw3H
W5JMQsQ//mL1pNN1yhuswdnGWROKWmcSb/bs9NJGgVekMsNAHBWL4IE725uO7/176nMoOeEpPTfm
p6i48Vn3h5xh4koVU0XapqRA1AuBFpNoyMRXGIeAHC8rDvMmjxKYmVD1jWDG0lq1BlZhAM1i2BDw
CbtbWBpeARAjc1uHh08Z+pj7nZ54Cm+FcXpf5A7b0rKI1FEykCAmAsD4jb7yYmxqrpl2pV38o6Sx
7dxwa3Tq2vqcz57L8vTcFCt0PpgSDQVvNN8orf7SMeE7gwzNoeEK8UGnTBr/77KnoElvM73DAZy6
aExl8h1AuiD3eNGGcMLSEhurcgsUgzxKW80iUCW2pfesrJiQPVfS3AkxIq02RbLyTZ3Ftg6LqP6T
e9C+6s+AFCeQjc57tdFyJ2Yhji6GdlndoDCVAT5f17YOrLW1m3UIKMRaTgV7qy3KklAbePS47Xzp
T/aHSsCge4IPviId6zfw963qoJVpMQPNAcsTuvcklKfm9egoJKJbFBnOb0ItEA9TNYoZ8HwhFbMx
cawvu4XJ5cjoPs5LuvjEMS0h1S3xEVedlYIDJ7gMIRpvV+EtOvkqwKu7jLKuDSU4xQ6ZwcHPP9gn
1FrrJJM5yfFQFzSfbVxY4ClMWs1VxSll1ANX/qh6ZUSRaiaGkBVWl73g4lRD5Ca2Pcx7LP1c0X6/
QYuByPFcN5W5FFcg2k+GXXmF7WdigSrNUuWzuL+GcP7p0RGAk5lQx1rE6P5N8RtvB96qVjLSrG5j
+g0j4ZNm90ihu7ZybvQCbfiS17dunlo+J1Sj43QN1sEzVot/ib/KS27vnXQHPO24zcfukdZEpGPS
tO3E9BkCJDq0TgcyicpW6OJG8LiGWnnuc2sF7MUFvEUbYd7xUN8LvNgNmbbj315CHrayvOUPBsV6
BY/cWtJOlIOCPRTXeYBzv+OwURsAunCFtcmudyguPUqPlCR4SJzFa6mGLIulECcyZRZG1t2WLXJL
zdkwjpVqkbEqmsFl5f1xeCZWRUTt2+FvgNaxljJ/pngtf924zzUGZErQx+CVvSqIsWtmN2Q4Ggwm
YcOBneSGZitQTVeQWqYLEUhnHsBXUVvPT+nVoRov5AkAHO1xdV/h9P5pSP+uyT+KC89yZwr2Qo2I
XAq+/8/8VBYJDzdjxR0QkWhBkkZxhG043clgLyblIIYpyLIOaguw4FP3OL696O0rJflcUx2W4J7O
Qm2qiiGhNB29+MF39bqB6aKOsVfqboSTNgYSDfh00famc1Vx9FsJ7aL0HZR343Da184T8LKow+Ik
iL1qlAbDL389/w4pzPxaKzz2CjzduW/xHiXzRUob5aWlB20xySxA3R3sTe/OcdHaki9G8iqEGmf8
76+mm9aBwIAaeSXxPbX0jCibmZ/Ix8LQz8NtUjxUz2pIlEG/9BZ9AZ6MQIzaQVwBBpTKzPOpGl35
EqgP3OksBG/cu/yo9w0XKC38CL4YIdydVGPdyUeOaYH21H0skOBbhpGAbHiF24jmsq9GJ9snHZ0m
R8y+M1syn7t0825m2T2ckLiMU9Kv17tSKyOTpgstkCKf9TleO1N7kcPm63oMsVJ7skjsyKC+soiu
LjJcDe4nbVd0O5vfGjzeL9IdDVF3FIfvWXVPdfn+NwQtSJdNt/pZiljX4bmJQ776a9G8xazvJKUg
6p8NXhooYiAGT30RrTdwBfgECUsekSxMexrMmevOKTwtlez5LkpfckOTMXGbyX6/2C7Yf/5CjtRR
ihTLQMH6nAK65EfQPVRfbdFnfq/YsrmMTlwcZbhOIQ7YrmeeU+SFCqWPas61w8WIPMG67ajWpgm5
7j+ReOU03y6lEZZkC3ZkiVaBkakvAJ7aAmbv7jcNkLvocsPrj5A0PWkfp2GPpPHTmg421zmGTQKN
5NWEpmJMSBhVrDqYzvqMjDjytUABxxcP2+h5MLKMXJCIOmaV8SnsDK4g1FiFZHW76kz50J9HgEfH
/qFKbJb/+27geP5KM3AbE9hT0ddgubo5y1Y/XSBslCCom180PeVM2lyMwKsswjALNsBFVYM8M866
+QP5hqHBm1PZG7y7B2poJ4uMLk40kq0NDfyhmhYUeWlGvONbi9pC+7TWVCB+a1MGPn//3RKZtzHH
LLEaO78HtMVioKv9FRPasVZjkqFsI/yZbVYxn03iWKoxZSZDRQLwbonUPaK06xi63OeaMxrkvmq5
MJgnsNKIp11R3yjgFSKFqkotk4wY9+C0yjlScj2v1eRAF5Upv2QJ4l7Gn5MRTyeS1D1719aGcbxO
TkAcCzS2n7pVJTk4JRKTxrkUe863JQqWR0JcBIS9Jb1Myewh4e79K9mHwa0FUElNdlixBn0uoVqz
0hBTHqRB6Fnf6Op+C4oXy2TQAORQxNfW8GrW76oTS/Fty8Xf/YeYoVCTJz3oizc/CVsNZ8tkCD/K
+zR9bxqcExUibz3NsJMAzpcLANTN3ZQ8yijqj2LL/Rw86jKcXV/hXfZcyt9r4YgX7LUyfTX+Nj+Q
d32PtDLoWAWf0e+HV+M+hpyxG3eC/Ki7L5mOL9sZ0+kp8molWz3wQgYu6y0rsHYVXIEj+mwwvWoj
6ZV57mCzNZiOEu9cTJTnXyNTyu665h+NMRxg157hjjrRyeAdvjKfeXed5blMyQhPi44sLZtvnM+v
Xa9d9f3MHyrkvdzahuTJL8AwO0zDWZt1Ai5u199as2Awbzx2+GsqF1q52KtphD95P3PLTDUaxXXV
BI3+0+YYbAGkOWSy4XtZVjBiA8QNXG12zEamk2cQzCthe/45h1xh/K1iWqUVv6xIqdQpl9umWEhS
BKnRnb4KewTbM1oGTuREvE1195cP4t840w45TzMztMbt3pv13eNkOSHn4mokW31gVLvZd+ugMtgZ
ISIpCdorzJvzQMhNAXl/mdU4578dZLGpJeyRCkGQ2b2DF4E6Jc0HNvWRVnxr+cQlfQOW6nN3OGkR
lGjP2E0iIJCE3C61KiucZ1s8TewiPs6u3aVyYrreH+lRgPAQuKU5/IzzyYqzspFbPGEiPryVBxNF
4UD5R9TB2nbWzo0BHSolBaD86ksQL1X5ZGHP6f7ARRB+efat0nDtVHsuWmIEIsnxikkjsspdBDIv
po4r3FY4Vw4XhTDONLv8zHefgPEpl8+Re/37lVT/jETjcllDcmUZ95dednwDKi4zmdfrIVVygyYx
ni5QwqMFQVIB+MnleOKRTy2PHS9E6+W8l/GoTupQuuEafvnrpXqy0poTRnYXygZ+9tYO0WtL9l7k
0ZoRvSZwydM3SOa7QdhlFNzLIlMVGVRg0Aan+Lw0j8xMGOBLAgIIubA46K8eht4PCxOCkxefK1Tt
0VjzOHbAdQ36XKPU3Tmdt/y+PQnd/6xJ1OnjzwdHEpoG0ypx+Rkr5RPHyTpQTG2f8iRm+tHdUSH6
A8mULbEwZf69jKfgohoq4xk0kCSez2QC4smYz6mXf7SSSX9tLpBm5rO7UEX0/dae+Zf5RKBovKPG
isv1t+D58TVV+kRCvYhw80OH972Lti6H8Kg+8I6WWhkN2X5p/0fLFDeSr7va4KdpiH/8WvCI+Qn8
ngIByH7mF0jhB+yXLTA9z3tCRiWjt7KREaSN1DH5j4DK4+53gkbpgZmv5AtPVHc0CdrgODb2ztkX
5vixEQQGFVBdg6BSOTVs3I2j2oFEfnKvS/94G43GMJbXVpV7vEZgHnj5/wrPT8cor+8BZHFDCkP1
HKeyicBB/gYVHgLsmZ+Fenh1JtMvnYtXYwE9D0Ks23lS2cDWHTQuk8xtHwZBvSpOg32l2w1Q6TfZ
NEYY7zFjyq6atpa4yCNB+yVocVLsvRyhsAKqyGUpGtFqUMFxxJQx88EURYXP6DgEltGdAWlrPpTk
qVq7euOA86Ga3QdrzxUg8w8+nzIM/B5eemgJbvzoa09FnYpM9+8PTbIOOsHowk1LBf/HqFBZ3uAB
bzCU86OBHk542evNPXt3TiYqjqPlt6wPkD6hGwVx1DBlCp2B9nMUcRf8QAq88lfajjnj8zZGnBt3
dhBop05GisKwxNNq3CEdtd5J8+zUd9M6biBZBXwKuC9lTLoWAlZsEZinBcu0Jws+a8oIRq7f/IYX
s+G7TF1olqo/SobYSObjy8/Lt9TvvTBC1eWRS8Fg7yZp1k1IJtL8+Sqhghll7rvtCDxQxa5gT9t+
T+3sPWJAXs0HJnP5x2wXvLO0/fhMRA2bZFzf0l8V7Lg1IEamJ/YyavEtPpa6UG9/74D4tacB4vY1
brZvNQLzRyaJ5lA8x6v+GgdTnBhaTThJHVAv2BXqX7gCNQQ9BIA+O2mSAxaCHBo3IQW+TtM+IYyq
3Etv+Oud8j9Mmt/9KlLQkBzX9GWav2XnQIr+RRels0ikbw6KDXnabn0EYDVTnSXBCZ2wCZLEjH8l
Ucl136zyuPPNkSoEyud3QUB0jcm6H7wfLN1fui+JcBiRHj7Siz7uWqIcf7RLGL++HsIPDCBT+2Pe
MmmX/WRfIQCsqkS0Us8DHB0luG3V/w1dQkHSvcJc25c29W0vJ9Y/xS9orQOQxW8BPX3dAKYGXTNa
G1XIzx+L8TZYh6dBoMeKPyuiceMAYJAh72hRaWr4ZZKOtiKFxdu2WnohgtJn6LQgZUVidCAo84yJ
UzmX3aP4LVV6D3sLQSsos1GJ8P2eKJVvE8EzRIS18eXgz7VAXeSXy22lQPnosTE79GcJWBBoeEhv
1z3TyVm8JgqA91+YhWe3dfAoUTdHmMVQPlBGv/UrC/6IweE8krfwrJ0i1+yNKzXBGOKo035ptg6i
jzWX65DWo8r8Ci3rGo5n4qdQu0AK+8tk/F07mVhi3awbtI1Siw807MXSO7EW94ZzM6XelvLs1ffC
0A6Q1vPllgVmhAHznbxl7uOTUYS3oW2U+QttWD3JRhT3cp/Z6R2LS5vttLpMqwNT/UgoeUC2cohD
fm6kfrOtYURtsXIEmD1yTD2uJtAzA3MEO9mjmSWx5sIkhPoKLUpL/k9ExENGXmWvZaWWFqlxKVrS
FOPRaHTLrcdaD8XmrXK17eH2wRul79Dwz+QT1K+ivtrKyDuI9/4Ya8pc785qgjFv0RKf2coTqQJx
WwkY3f+fMt5s/RSIL9DwUnPJ4Ka2KGuKE05txPIxywADtqWzdHXmrRqWpmkXkrsZSd5QIaXaTZPE
aQ0q7HAzdMndhSZUveKUOYLjFJeDU5VmsJUhxPBIJcx38sK28fPcGz5TrAaUHy4tUtqiRDN9noZI
edXpkckU9QCwq9pahiD99ileJ5NUJLaaPSFl01Zpb9mObaqfwPSC3quYiFnEuPc3AzGKS2txvrBY
+OCgGl7cmKqxwhGgyMKM11UMW4O7kEvyYpZWh/HMbtt8EpZpG+5cxoIhfCBkykokxXRnycQ7vjSi
e2oSX0mXAbAdv2Yn6L8qBd26yOqHa6fPWt6/MqFth9jSPte/qG8mcbN3yyly1m+FuXmAYHUgSM69
WWX9vKDBTkbL4tKysvKqzraWN+VT/nXeYrZM7OsSdJLy+Q9RwkxCXzE1qLar2KeRz6ostdNBi7qC
wn+bSr6VoFd2XiM9BA2glKP7TTm1L6A2Z98N0kDB6El5b1FA9s5FjW8jDkfjedMoPonsIlUMXMqR
H36UK/9o7ENfYvy8nsHU3sw/g7hWJM8d/tmviAOIGSxYD4y6kgytE343Op1jGY4KDM1jjrk4DvOz
0TGH4elMaLOre8Wcqn029WDWWhBXBdeO3ysZHLS+RlO5GgbFzYYNjl+8UYJopaaXd8xyH/T72BYl
SP7dfZ58QhAybNlFOMlnWZUhba4bkeMkpZokyJXFtoOWQDoxkJOREy0HQc/PAI5UQntVTRFdc0LR
Dri9pTFdUDVfIw0mIHhRNtbibxZfsPACLnER3szoGZErYXx+dosjmgsCOCVPvQAf1MmkoLMNMluC
nJkrkIJKz0qD/qAIHD8umBabyBTY4l0ysYGiUXEWe+OAdxgWIHzWi2GQvlyK7QMunCAJZiKCu+yx
PRuFFUmv7QyJ7nV2U6G0XwPcpu/nG9iNFoECw4xjcjYGhKknpIaazDSn+MiIVcRZSQ8DM+5xeFeK
8nKt2gIvwMhIJpJISZej7kyzWGe4A/gaFUJ0bZXx2qg2hd4qZv37yNqYWw6W0Ke0YN4EuSmfc67P
n5dbeLOAb9krgOWp4x5s8bE4E0JcmqN13pJ1+GZQVgND2yzuyFZ0H0OgNnk0pAwP5fiSEnrjRBkP
qEup6I6/wSvd8w6ZQaspvV0M3EUq8/TwAszaCtKUp2jMfnICJSOcNMVAE1d6Qs92xTr69IpAjo39
m630N/xKzzaLauDTolBEeMLmkQ/L2KRQciMQyEN/MYqUahMP2M0VK29J6zj92+WQSS6mO6/BThgE
QYBiFOh4BLQwml3B4Hq9Dj1l/lhR3xEoFmjdJa9D5tfI3UwDobiLbPVcjjwR4Dpbm/wxea28LvaP
Y/UdcjWPZCbWta4N0TrgTYf23MH8atoT7wsuU1R3OEoqwGkL+CD9xZ5H7sT62CsU+fI4voJG4baS
PetUC6qLVBJQU3GrJgEhKNrmWmdCx2Iv8O0iZw2NTODqiiF4ctXcvhuC11DTCeaol2qn6lIjCWuZ
1pNck6NYCjbcwaSlG4oqb6A5TYzTJHBGuTqgLfSOVbSvnAgAo/LHi435izxAOgXbZZ7SE2c+qyQi
hGLgu0VFaRGt+I+bu3qhu29xhzt2DwN9ipFt3KjUk0E9nAysAfUuJz/lk8Tcjz2rQAKCy/QPl15A
UtN7AcvDfEuGu0uZsjgQb6PmmphDYPVkHnD5TsRI5xxigNHGNzgVIJ5uwHPyuF1T7sYrX3mhTZM2
U3VJgnZW/oFrP2vyLkaX4AWM6NKpxTBtTcpAHs+HfHAukjBYJYnB/BQQsbf67zMICxC39QJGvTBD
uvQIoOWs9rcfA5s2y7Mcw4g8Xn5MiJqTajK/9F6BIR6MFZePztvWVzgCpFigLWp1iUEsCAseZwcF
60hON+ECqC1dDvrdsli1mMnCdNgre2udw0BQXHN29dx52TJTLc/NSOUG0n1O72+FVZiJ6u5FPyKb
JmZUUNGa5td8MLBcAe/R9ShpCn4nHRBjq02bdlBuWCC4s7QyTUC7900HTgMMNNamOYXLQpi0DGRg
HpONdJYa3dfGkmTnUkke0KhjiEjrV0GPM1kz32wyF1KYiRSmKPRhbJWOS1zTFbV/m/LAhtJUj03m
QtXLRplhLEGpRdVmbS2zsT2eu5IFDon0NJb4YrUoiuQijJ/nYg9A9pS7nzMFVLJQJmqDaJIGKkXs
PG9d9eIQJipqKPZYqsr3tmDRjc6YBWxpjDMu+lC+u7yM5a0Fu0Yg6lGxHaB6uoFHd8hM3pfJoWmM
BdQsk2JJSQz+GSOjx6TAu7+KKUPJbac+JpvWVigcvgV1zMrTJhLdd1hnH2WIYGnnxjS2ECixLyQj
MKfUPOLVEA+titZ+p6jAvDWVjOtfT22HsIvy/Txk17x+xxrX15V28WySj6TAeaUC6M/+boTtpry+
nIZTnXoGheKLRRfr5C+7iMdItAt2tl7V3fPNvNiimXr3tXS7afpFQmXU/W4G8gmtk8rYpFXDYgl6
8JMpfZu78vl+EnKRSiB3DB+1rB5iM3C0AYAWf2V2wKcpeA7cBrprE5YDC/af+ehgTb49H2114MEH
Aq+OqPbnyIMajXrK72LgfcqasvozSk3tCym+eTmSm/vOlS7l7/Sclq+h8BH+E1RcX1a3+q03XUlg
7sr9UtPLhKE8ecnxRA8jyqA2enXdrlMUgJlEP9u6VwiGPXces94gCjhvwEqOSfm0G2tyI4uj0t4C
rPI4CIDfua7H+3w8rk3M+T2hNb8fz5wvESQs7CcyUUrZ6b8mizUlvmBzR9r+oGdDIl8nnuAlzeQ9
TtdlrxE+2FaASspcRoNF7zJ0F+Bmi1+MVSIIgWhGmOUt2QS/RczpgjlK0CYjhq8t1UWKZn8jxLM2
cvxStUjPiXZIkqfRaGOhB0XqqsQo/5Rmz9cWjh9On1gryx500xnCtozVk4jNKvTOLAXR4PEG3ppl
VHpb9O9y2AtZ1pod7yphSZDIq2z4eJDPnO8o5rdppwi7Y8Ryggp9kIF2vw69P0ePi0DD47QAiarq
4vRE0QarYpCS0d1jEWIJfZ5DzClOHINjO922AlqeNbDAbV9leQY96Hc7vv2ccUMJyhYvk68E8M5B
ZRaYTv3H+dt+LS+kTe88lStd95TULJuqXd+AbmjCcIqj28MJe7igqSnd+747Ycf55J8XlCjZfXX2
oEaReY23rwDogwU2rHiXSi36k9Wc5Ysg7Hyx/JDp94qopbFdbcdDBzp4uXA0VyhMoEpbTfXOCdo9
BdiBquxYRd9R8JHthoQwB06uyjbZy5FZzA0VPiB+3jeSqDeFCAXbWy6UoHZ1k8jlZWzvcH4AIp8R
3/41WH1T1QIijQs1Zx/s9bjasfHlOYV8vv9US/JXB87aYNPfKYuv9QFy24ZWrBQ7e2Yq/Rda9C4N
JniOSsdaz8Doo7G8GF2qiyeOQmk4lXkYQY9T+t7E+UHKVYw/v2WspkcqE/Dv4XuPSSK0VMb5+YYg
c5mCv7mB826yoGKTOSXEeCCKMNCyR9kegVELa1N4SsyJwk3TT78V6tDInCYqBU2PTCDmILyUoKdp
K3sKfCtD1PLZFBZ6rRJ9iLO1BsoS2uQSEyc3NjCvjCrcfVjTjR64xnZYrTSWoH8sskEkRplvlTV9
a9hCbPOMvZzMUdmUU5/UDBpJP0djA0H9hXdxEybKN92Jx1jBQ8fCdk7IP8DYJYHHPzimDdagLPV8
Rjd3q/Ez2oYrGmTx/it11EghLxSh8gGfeuQDaU/l2naz9GRUJfdvBBR60r+pw19gnrJhm6E0g924
49wPyQTThJLnbgf+/vWn1VWh8YvdA25p1+4oZFHfaAmKM7SdDa6VQZLns7vQbuHZI94AKJv1VpBn
fIzVo/yXNBRMdd46+ThqjgvciTXdzMMZaxZLVSUcRwninmgLGSfq4vJKsQaE1iJvY4YiItLw4HGo
OUXjOkotsv2tIZfBdSx5VrkW1um84Ejj2NljS+cokio7g23CLfCr/5roswhMsLFNt48XxlXdAg4m
2H6wuq53rQnvQwz1G+9ZFezFfSYd57VZ9MO8Jdkm3BLsUE0jKkZsiYHu+oovT91BXJKgyk8YmjDF
ewnmQ2OAyy1QbYlyl63TKIvyN5rgBsDmgY5c9IuF0QDYEq2BaHVyl3Ubz0EU2jyZ/2lS+OM87+8x
7d6M78HgO4hkr0Js4Upx3agVrMVQyG5Jv9L5UF4toaukZcpmGVlc9tpY+8PM+cPE4pvFmedtT77g
iCaT6qYkdxU66DrexZBoqrwgfeqPUIA4l0Nd9UBVBUx1MxVSSNZ5e3+joTK1PCp9KcOnRfFbF3Nr
IHt1794lnJx0lI4X3/aAVjxgOWwUU+PfLibwR36M0zAG9Mrhu0c7l0NECwLOQYVY61BAOrqeXd4k
HdioPoLWKVi4RJoVrSaIgwQxYjZ+WR/aqAwbhW3II589X2sk3yFltiExBn6BQk4oJyZhnK22soPO
d/u54rvQ7fZLMK6NYlOcuA3I50+H8yNvPzz+frw7DgL3uvSGrPXLv7WHaz9a0FaRImfqA9TE0/na
+dXgYuyiUs6X6E+68Huiq1IZ4j74dfhPLC/xLKS1QqgFltXfpaNdeIghByrML32z8ordZVwEvlWD
IMokEbfvCu/o3QQWZfzH1xxjy/j/L7zY1O76KbYkbvU9IrWlQ9b/8CWYWzcKZfmfgHKjJJyOSwX8
5ciDnqDyHsyAI9fdHyOu0mhkCMViupFF9zu2PLUafca4jW9bCcJEH+A7bMWo3Ix7d7d+re0o1xJ3
LNAzusnk7mXn+YIjsBuX6OjKYUOKY9pyg99HaW75/wTZ8KtJTrxnnQgXlJkRNip9axJlsHEH7ITY
MHvipFuv1xMDKJS8Uzd2m/Bv3s/Pq5fKThUys0qosZ+sIRUdlo9MMXt+3aG1gRizZLOdw4Ay3NDY
vi6h+3A3VmO8lLVH/Ws37IxAy5xQcXnBwDLSbw2u4LpdJm9y6NCBZXR4VfMkNmguHUwced2TRsAi
ERHo5qC0yZteiXnDZMACBCSO9BN45UlIuZ2+MZONzqI1oXc+80gFeSBaABcx4pF1JlBzJS2DSBlO
6OQO3+WA4r6w/OAX+GR4W5eEg/5mYHV5kioY1gAj4UG/+RrkKB+5B1c7XRlzVC8zz5YQXFqQKrWD
cesCE2MCzx5PLS0z6/pxNW1S1XxD8u6UX7mKJDF9RVgS8X9OWwhcRe8z2L2Am0Pj4cAuYyPQQZjD
zORUB+U5BFwphWGLIuj+Ac5PPdx5r0oEly4fVp6u0IJvIEpHW5oElsK88Gcc0oVGDeMjbeeXuFrN
tF6tPJshzj5PRZIHQfgPrqWADLklryIz3JcoFXlMCsrV5qRIQLNZSj5xASD/D1TDwtGriCnOdYns
R5AmPWLm3sc3YnFpGNfIBxQB0FpFvEkN32kwiFzm3av5zV5i28RtkGvWX9X8bpE81Kuea12Hjlj6
rMOy2BFWngnsKeauEPaJEyGmNPdaC6Vq00wAVYnr+sOjWGWSPH3wT/D8j56ksPA0h9r8nuzXrPM9
lEfEHDY5pf1e+MEXlFj3eFPBvi+9G18+zZjvKL0OEd8rq/Yc7MLt/J9at4xA3rxALVZfoQWA5MNT
LmZqCPr1QzFydlInN8mxKXdk5bZV06T9vW4XqjCbja+tx1WLYI8TRKLpUqaWtKIYuYR2qfPXYcA3
LmKjT4yr8EcccfewS6M8oe3dQix2Zm/huZgXlcCfzdGtygoRr8rNOTfYL7cafMff4VoLwi729PtD
bN2dRbionzqKQ/UWUhI+2cvPjIIib06IcJsVx/yZ+pQvHZpO1JNEv61tpjHBg10SHaLr5qji6A4R
9WjAvuc4nmlksB5AfJoN+jR4A6I3vYElbQNmrUYbTMlsWCtp7UyozNgwY1RTV+voAAusmUQVD66B
LEmF+3QOPzyFpGf15rMwpwaKfQD8GuUaWWTioNFodEX9fHokWGLypqRM0vtB1vnmKGdiYghCV/xL
ZQzWB6KDd2SvnuiWZvSfPL8ZssRtUagayjxwubDnxS5tw6HL70lWI7pGe3nJ6X7dQBzyuXWD3Ybv
NQibV9Xi2r3nda9mfYGNVp/zA9UdqOKvJnMK1ExUra06EEP7aZb9kH5uAFo2bEDYovvkCuIlAFrS
cD42kqVwgvPtrbu4qsSs2atX7fWR8rMiiSkfvFRLVjW61W5+WZkl96FFmmYE+r/b5lLUdT32nUHE
7mUbliCqXCQyG/Y7Zby/H8JCZI8HEQ3eDhy+kVdPZe7fdUk20zOOLuAS6nObqO2N5XAu5FXtNiSt
PUe929gvnLMB1aBUcggVm0pSDnrWwX0B2Tc5yTKwj895usZpVf5yk3vUXkEU7nC3umbqrUhzdzh+
fkhBuC3rN/G8hXoJ7t/Kj7MCo0cfeZZwlH9uPAd4gFxUZWi1Fs8iaDnC1xPApYPvUanKrWFcJLGb
XOmUkxO9+LP/7433IbhpVBNpNk0Vwcjn6huDnaY6TF+Vnr6x41PUDVDQL+wsQXs8zfZu7M3QE6Ob
VXl2N5cysYntsQaKd8yupQcslpDEs4eC4pp6czbvhUhYKRg9shBlDO9XW2XsmVeeZk6G4GOtLnnb
lbK0n0tLeezDGXudaCUsfzBpF0aEqt6FD7Mj6rPkhC3iZEnnIQqIi3KkXX14aZZnW26xazKKjmBH
hbnALLOTcFH/B0ss5aePAu7VCyvAquhbrrdh3FQgzF+Ss11XBTIeUkumZ/+C72QH5wHqopkT+URc
4KR1Jrg9TToezUdH7kTKWDM6cK1RU0S/lVqrGfogH088tHISr+Ch5Fc008UNHGuI0Z8GmjScrMMz
HEOG8mZ5WWH+/sevChxHDhTzfpWjBw8MLRwbc2I8ZsBbQYIbcgHYQI/y4H92gyv81KxnZZl1qiSm
EU6EShUg3o4RbjnGRhy+5RnlAJnmMPT7aNlReKijvbYcTpAZksluJwQUNMReH4nuRTK7BM9ijFPa
kYJeb5UA+djtMuOO2OKvcPDuy4wLqCFW7oGuZsmxuOFkpddIBZXUAGRhIbPPUVxNg+U4T4G7m7Dr
sfnLfrkzjlRHkK4qDi/aQ9fmoKltjNRo/tepdXAgObr0uEMRioSPd/8tOnD9HSn7m3e67Qdk9toV
dpBLvo5tal1lTPjUIcueIKXpCcVMcIFKjVXLjmFG5e/iFk4CTAoI/dGljxGotw8IDC18FeF44tM/
QS72uetlH/TP/5deVZ+7mMmRKtFg3iI1prnABPGLvDrTT/b0Rw7zrUPxJQ2nG3mCGV1yLn7IWRw1
3d5CV1TSg8/BJt9kizqeq2SUiaLtIFuRTk0OJMviajmbn4EMKadS9I5gqxiyz/+YjHASl2WGRDc4
8vzVeZzr/74Jr13GOkfqCVOR2V0e21h+WE9SSq5dMo+t33f547vaZ7LNvUpHG64PNEiFhKYf3kUE
/JKcpr3YSTNTfalzKIHhSPMeNEYgYgqYZSfg34wNUBhU5CcU2qfC4sq6ihNQ5BAbjFPo0TQ3BDuv
tsga1dF1BLoFKmsYQC1jH92IC7eJ4Ht8yoraj7UcqXPUWBrYvCAT9EC8d1WIxVFCsy7A8ZtpaRHB
wXnjuW7GQm3M9UGdzlbXSNAUTFd7drDmle28F3lAHWsTLVixYjJtB2OdGZQGFSfCkUBRo2hLFCtT
re1h9idAgEJCl2s9NtwwYdpNWYx/ITi2H44gMeJ7fIv65wlQyGrNCrHWXQYKt9QndD1AOmh9vI2z
FFs8/HmFsCwXwDOK2P/yVDLfPkQUBh2CRsQShLNZ5FSXTV9ap38eFRcfgpFbcXheQQ4P/NqDuRhW
ii1BJdXPMuD/CrwCpefnOkKX9ns7Hmxi8rSAvV5Xu4sBi+/oxQ/eYKkal0DypMIlFN756brXwT7L
1kmED62GXshaqwG9x0tKz1EdvJrxS4nkUH9FZ9/+hAdBBW5sW6tvjDEXeWcS+5lbx1juSbEMw4eG
O8KmH5Lyxhrd96UtwU2ECcGDD2ItZddPOOjO1J5bneO/k56QL/rD8SJINeWJ+6ag55cEN31u3PEP
pzPagtg8OmiLViCvpQOtiSuv057NWjXlfR4HxwSs4/3nvcO29o6pHdnYDP7AJoN50/y+8X9ANJGL
lTLJvDhE0djUD9I0uZLY/LQMZUif2xY3I39MBKZFlEIfJCNiyOYwl54913gIsGELbYrkP6wvEUoj
x0Y0qpAnHvCWOYXUxR14rsPKbH8FFCtKY2TgCSuW6Uh6F4F/px62bu82CJ15SBTZg+L4eWagczoQ
qbbJjyzTIyPfVNnrvuInuZFQYgJahdjSxkaTTxu+LgE6hk4dIeftBKN4fRtPuheT+r5hQ6zpGp1D
UHytUcgx7iKzJUpAg6iOZCPGQWYFAJilnCDzqWp8M1QJJv6LnrXnKF6nlhllIl+hKiwR6zfeDPzY
appwMl1RGYCvRsewg3JHNfXNTJmZZTL4IvguSED7S9OXFKGSSv69SuiDED8WXlhaWma4YQ9Lipa9
qUU2TWvd2F3HYyjBua5z53nb4dirOz7JdvWOnDHXKS5/xjbLqFUHXZaNMw+1GCYMtXZkte/KyXCR
nNr16wT3W6V96JmQoHckWIEEHkd0lu6UzguA30TpabqbLqVBxHSG5dVO89RUABSFdte8o4RkzObo
kYWtGLre+1NDF/nPTMQCTSH8G81vl0upKaGWfaa6BRstNsoCyvOc2BFwnUKPxZrXmeTqkR+HRPQ8
4rJKR84o9AFJXapqhoiVmxH2Os5rWXxOkcx/6t0Vp7eOJ11TWdJy+K+kloerp557C2WuazHyIKtB
SP4rDDQPt+apTzrj0qDQPAqHwjyOI6GiGaS29yNKtY9S3HuWRD3EuGo0bbI8NDOAf2ixxXqrs7BJ
aN4iNGS5myDyy6gYlHXwIjdcMqWQz7PIIFDU/WDNzUIs09rtroM3KhRO+UnIjM1z4IrXNNXZh0XV
uAU913Ql/c2ttqajFffYMftn/u4C2us9ZEFRIWwgGo3x6ClOAA1UdgyJc5eABKafnWwi02kJ8+DR
cD+2QMXq22e47gS1h3MjtxGpnr17KXOIETKwQtspj8Ed7xmXN/PyTaI/iTHeHcyLwq2CA/JgzKrI
p5szlyu6mzq5fQIqzlGYgngwwYMXlPEJBKY1hVi49NvNMiKz9mpjK3fwfcOAKjbiqj3aXH18yaJx
/gpGK8Wkbp/rKWkThO4KTVxrJkPKFq7TQ01aZwGi7EHhhgrdXJk+F1G+Jefyt9CZruTicAKrNHg7
5UBB8s3hssLPQ8meIM9hHurW+95viNIVPF+Si79FJidEpxXE8DhBeF5OsmrABQaFeZjomB9KmUZ8
2mLcMn9GAwzR1jju3Y9gckDrSVGj3cNd7uFRdhZ+j6Fz79x5RP0S6uJLpxvKFnqg9xBGVgs3kbd3
PsCI7AMen8WS8LTvKSEtYFN4qc7rKz63NFP6NgyadiEHGUROCjbJpgR0E8ImAhUtRXvYJd19G8qq
zCMB4vtO1NMIo/bkgnlhCLy2UpOlfPv4a9T+6s/dom+/Mu7AQzsALJIxJW7CL808WsbzQPZm2boO
jmII4vxM6z+6ce6yKF+LtwY4kUNkI/p0s1llj9tiBV5NvLndV5dHDVj0UhLaOY+35SVabKHkFMPT
vGOsMlr3zl4GHzKD9A0e2eL5kY7NhK58lZUWDSXzipCWcJOqOrEvhEX63+JBNdVvMD08PLyXXjRI
ksU+IqWJY4458YwvoclsT6htWIBlC4LqWow5h/Y4or9ERp4FOEUQr7i0au2tGBwkgSPmopvzvO9L
WcFN6W36vD/isQbf7wO4ivn9vIxZxUmEQ+aB1VfSuzQ7SnwCEu7JVQ79cfF2jFTjuX6cUGibfqX0
ug8tLgTnPb4oKPlAHYAyxWoANJaVnYqUeVAwSoBtrQCrShucSi/9fvP4lWl0lIWAno19+J0jXAAR
Orc9HOLujvLHTKJ2sXF7ucfe6IxY2OPa/8W71BUq/H09SitkHoGxRn8OgapIPZsZX1ICZh9Jssr3
8Rw+afM86/ewKvhGSZp6anr6SRe7BdVD1cezijcMP4bI6s4T5WK4re0duL/ZVjiaBmr1Zzk8+XVX
0I9YimGmiRclnPNOMbYzmiNQtoRL89s5yQ62bqEPy/MZ+2rKPjeS+O7dQyNF6DZb5XMNREOP1UX2
PeFwPaRwV/XD26Z6ZQHGPdpYbB8iAiygML5qasw1Yk8Ppp9IRK+NJFxQTrf6kX59z0CicR75qwYe
+84Lq4g7feQ0Sh1xrncRgH1iFTFMRWHg8PzdfPIspuAE27R9HokjhaR8w4wDUjCUxTflEiGZWWRu
8VKYIYEey9yEAxirGoN38TGCsJf0HpVWHMA3Dlt3hEpR2fdNWtwa9NUgkq0W2Dw96nsckyk6hADx
rpt/Swu9KZmvRC87h5ZU5cC9B3DMK0ATOjFLE1wUePBmnO0qgVxU8QQJJq1kGVDuMCSpdD3wtQIj
dfs8RSs07Wk0DbDsmngwGwp9PlwwmwwchMAE9cRnikITDgjb6q5McctEf03dlagr5oXfUhd4uGd3
unfnWJ9p820ekfXlY2RM7gViuqhkcojdVHfvEJxq16h187wm3ySv39gagDVCCXwOMiSYqu+25Y2p
v0a5jGxo+ZXK+lqxgAWusoGF8cW3N76GDSvdIHmeeyqaYCQt39O+J9aSaIEBWUs5bceGtQp3Ufvz
4wRfHnwM10v2Yd9ZGtHaTDRZDMJvQyuE9Tg3EPGuV0ECWPDTgcYh7teQuJ1CUsl/128QLqZgeneF
rC4HQHvFM2IxwlFu8Zv0wnu5KFqYWYXjHhJBUaGfHVojoABryfv6wRrec1wwCGELvQe4BKXK3V7c
Qy4jARqR5xprxTmBg/yjBTKUIBS2rWLb8/pClVqVBPYtS9e6afVZSQ5PYQQ1av7ZF5fj2Fs40mxt
+GBsBNcN3A7qkUZjizw8Co8codmI60jo9VD/ZcNpaSAKjKkrHAqEK2aSgxmFxk3xSJWiEBaRXwkW
9DWDsgKcapPt+6bNP7x+ngtlwjzIne/6dYW0DovIlxFXgEcNgHlZHS+3YWAfsnRwH7mWkxqm9ImJ
b678E2ovTM3c0wHLM8eR9REeYFIInDxy3Zr9+TDDJxbZ8Cn2ZgHNYOOGh5oqj+zGJ5mYu8j09lul
hc9EW3vddhQi+iwgkd+xMrS/88maJhu0bIuVH8/xXUAngOlFaNaiGQPJmZrlDEgYWyaHnal4uLGy
iwiJy9erZHDdVxKLc1+IqObGt0f4hsHy5aG4Umk720/x9YjHOaU+nLShGn7Ws0bkh2Z+b3MsQyNE
t6DHKJGabzEXiDaTYzLm+htPP6tryABvTGDQO1pqD3iutcb6JV31vUTisDdFpo4EVMfTno/MI7Ww
uCd8/ZFE6YVwX+9rJH2+1sC3vbFcmMAS8qEuqFtUDwLqTc2nWbDuWkbSQ/7U5u5V9cL7HCS44KpN
nhJxFkLYxe6ZK+r1njgvGO17vzB+QcTiLJ2Weq41gTSZHpA0A/T9Y8M6o7woKYazewmOWyrqB5IJ
uQtHsqqcIOjXrFDXEsIAYHj8KypaAOhC1KhyVgz7Ff1INvEuIazDKMHW6CSXSVj7pVa5nMMcpG8B
neO2u6POEdyqC59j42bzHO/iiVIxjkIOqnB6CgNh+gBZdBe4DtZYD1g/Jc2JNDk4ntZET/R4mpS0
/I8furdLyDnUOY9afC2YkyqLNTf3Bb4Z40IyDLopZJzlttKZpXWdrmcEAUnfS7NGoZ2N6+oAJZWw
ivDVIMFwBd+YCVegDL1M7X02aTGL31r06UCBVwe890Z/IkXmPdsXlwpYyaZ4TW3wIPNLKUM8IYiI
Hfeqz8eTwzKNbxyqp1RR4k+rlKG9Rw6yXZIFzLET6aQUaQoti3pGruiEr9hZIJl703NFRVJeBUwT
CNf3C4SUppJ6zaD9pmrIowJ4OMkjQ0ab51QooV4mh1WFGvWwAq7Ca94hAtivtGsRyMi326F3zqNE
lomOEnhgSGK8wY2FMFt1ndKwu4ZIJaABJ8i4c7LtBJv3SR7OQOK9aKD5IH2fl9jrJXHVzwEnCt9P
cl8rHTmqdCMCzdG4hTShmKYlLKIsG+ITpmiJhEh8hTzu/hPg/BDplnlDbs9utTD619gTOWNvGe2Y
5kNkLjMifZqjTTHxwOWTKq60aknWthOEKIgWyVCy+oJCqAayhXjVxoYPROzSK7FnWlnFmvD4tPVo
s4FPqM7ceSHXUobnSwUvg1d4uMrrkzObR30dqCOulUmWoYO2PQzcQ7XhEjby6y9LtWcY4X5Nwho0
BkruPQUd4HNmBfAqigvRJ4qg0aydHrzjjoU9AA9wRVYtuqtmzIlEr4Aj9ZUE43lrZoBBCZ+3XMzP
LYADbN3udZ1fLvAgyLrO07jMgYcnUrUWBG6l0HgVyZ3+uPye6tFFi5karUQ6eGW3+inJ24AsM/u8
Teunlj7ZKbFlV2PEG/lMsINg6fqt8EXJw7eqZ+zbDxNi1B1rST0lzUFUN+gv6P+gCRsyoI05NsEf
8Nzb3Nt4zJsk6Ezw/vFzA4yLrWu8FNAI3FvGC8+OV6BIv9EM2Xwl/Gcz9hdB7JPxaemcgauVgwRa
AnIDU0QTb+KiAeVkhYR4blVPuVioO/o94FHOIFESjc4kuwq84o2Zu66ZnhRZ6M0Ogtq+attHD0Qg
VO4oRElVjCMTFuHNkO7tVBa2KxIWIhAZOaH9EGsvGIUINgN55QOjeenrHdCAyZr98LUDMOdT1/3k
2jM8ICS+v/IaeX5l/M5IioVDOerAUoqBMNlptryD9+oMUrTPGnQROUbqlgelFcJjzJg3RYRKWgp2
zW8SLLLZILmlOHs4QZhmNxogUjscPX8knLCN1PqxnTBQGfsc1X+WG4yFVjsiL2mrgiMgPJ9MhR93
guum9wSkYNR/YF5nbEudsSRqXJErdfBwARriuiy7xA/LHWVp3SXZEgygpGU2seGVH6Th3HxnHptJ
f3GWDULgBZsfs5KPGBmj8+lI3a4jfE13rDPsa6772O/UqP/r/HrdvcI258FZpJXSFHpOMMCoUHc8
FF04XPTz0R/x/BgoBDT+IYJm34LRDt0+28dtTlQ/8KwYvClbTu2SX3jtQHNyO2jv3fvABhH+p/+p
t1I3ugfLQln+0+aMAXZIO5vuJroAbT8U0XBneQ4RGf648I9GiIS6lxG0DqOciRtsNNFaHxZCYWoI
8cENXPgaoRxpv0sNA/FSjSndwz+2DZpibzHiOUDr9CqjzjE0sDvb4LIT5BhOF1QqKtn0kCtbqU9X
hJ26h6bk9rBTdirGgfMoNsAMsmVFGzBwB6TfJZuzxgxWli5hWnGlgPyiTu2C7X6bgOgdvzQPLK+y
quIq0DF7m7y2d4NKfE2SwBJevsiidWY9ggzq/P776CGg9MXXjPGQk2dKGS0A86zkp6UBIm4sAQrb
cB/mBo/udAd7KLMeB7IoT/1ig2+nWkbXOUddsCUEPypw2IeqQ/5mFXsKfUF5h1Z/YyW0GYGLQjNZ
AOjoBQHUfJojd1SMrN7hAGdGncjm1eK/VcJts+d9fJMtrBwGxS6DSyByltcLy+WmPRrMLwS2TSUr
xdVfvKf5yjPpD825Znc6CWeB+aqqCZnSSABem6ACyEw4fMmSXGuIxYrEttmX0OfzHE745G5zfKWs
BmDP3P0+y0RWijmSyJyVC73qyei970zs0J5WiW+AgBEDBXbzjsLpX+mPLj2pdSq+VggV3+FYBw3x
AZyAHd7VshGtTog86+8Vv7CF82ywtkmLN0qVT8KkxrIjOgGX1/6+2MXwXD0+BU4sz7XGQokcP+va
3Topq2+HAclihMba0br2W7LQPNqE/PMApUC9R3vOY68bJ6qHlokPLu4gnfZiLg1qbsmA0+SO6HjH
c/gK3+CcEhD9IgDJ4TMDAc2kBZ0ux7TssMuad52Vp7UOPv0A7WMgAeQS2xloMitV6n65Z4Egp+yg
/037ZC4Guo5Ie5znN1gXqXro/GJ48EE4oLtxet5BKGCXq9fbQDdnoNr7DvKpicSesoBp/k9clHQ2
Q39qAWJ5eM5lASjLVmr13gPyNaGhS2qD5+OJ31ElAragpw1oGqRh9HA/lXpPjeR56sBYnqG3A9+k
jz3ehkzEw47YAIx5aEp9RMWUJ/3DNY1yIrECSUtwp3RVvPnGhZBZeYbw+feyi+mOxcLk89It8jbU
aDOJlscO8Z7/eN9ZP2wqVNquXol/9J2y74q9uzE0guHjoAz3w6sOFaXb7EJUydSnkG8BSCSHVPGl
ruY7LrXQpFjy0ajTRRpbWhg36hww1mEyl7Ri00di97A9+/3gOi1C6xQjSphRoJtFPHg7KtkTzCil
R2M+lsxAbFRBQnsm4hS3EEC4YwIAiIAGXcNZuPUxwd3uMQHG+ZNir0bqpH2W7QXK+6zgpMioxLOG
9Cov0CTPtVrXnOnv42e8wRcdpnh8/LCYOCuZLdlJTLBF9Uj01UH31HestISHIapTMymAcxs7E0fW
t7XmfZQ5N4dLQmmtKkTl26PmeYrGU/SPf4nTT8pnsfuTQvfeUWK0Q0GQdwgaAQmqn0riqCKQskkZ
RIBdgjRzj2NOopoEyLXiinyX9Kz9GAJuvZV757YepX468SOmVtGH6HXkatlKwntk8OcTY5zhKFRa
/zFnfdjPOP7MHLECgKKWtM6dyWu5SR7leXNABiA5QU5ksLUr8t/W71AbtMdrfTQwXBfGANiz+aOF
ZPQjsrsgwipfhW5BX49jxPZbpMyVcyuT+RxuxRq3K+8LWJEId8pPUAT8dRC+8njU1lKc4TUovack
JzNwvmXa8OwNlgupVuBacwLQDTxEo8tFSyySkvycKMqq+2gH6DutAoHW9Mb9bkv3RVCsUY6JrDCE
g5T+bzSckALY9yQ9+Wdf5T8BayNP/3jEJqPiAQHJE5X4u9rExLt5qTT3q+cnVrVNUwZrLgAfWBtC
F78a49eaD2PGSZyOmqELZ1aptUTzj1dv9n5U947be2E2jC+4aFpx+m2w3lNCof8M+/IFOh5rPCFv
z22VibS7VRaC35roQ5eiXu55n/LKhRKHjDkiqXTO2KfcWQMaX9sEE3DDBEfyxJLE15bOnANIMUEm
HEnsQasvQNvRi9JhpRueJVI4PDecOAISpYNPcdh6ba3T5e4eU8KTMdezHACAfNwwDxc1fGtDZtca
4z2Lcbl5memoNrnM+7pfqLUqtvC9cOvp9t2lg100DUyoAvQNPj0o9QhcVKMpRMVFqbxkuRsXngR2
Yp4jsEZrdGLcX4VifD+ii0L+oQf2QnISnbVEhr0lUSvs9wLMhKG0F7mloU3Jfmf3FqJCsgKSl5FT
fxLyjW6CFh/tmrsmtU7vl9ZvDEY0XIcfs3Hu6z2QiKNxY6o+kuSQ6hlt1vPM0TGKU4l4ciRQKK59
5mQ1+XSHo56jb5YoQ7XaJe4WoEm8gtxPVhvsx6eSz9CnjBPH/DCQTZoouav7Gp+OMwK7pZSB1M+s
97acjnzZOfeqoz8qAcVllVoqZrO4N8inGWeFbYDW3oGoVtyiyvvtVwQ86almJvihqb4rqv8vJJ5E
u6FArbjwN+V0vrK2zMANlOKyjJReAbs1yARQTOvG6+1Ah4SBBiMJnuTF/f/lxt3scTYa7s7KwroK
TOnk+XaaVfdOI9nPQ6/UHHycR7NwuAbwvpTXUYf7R3POt+0Ab2mc2RBO1WnVLibLGdG928I0RJxc
Bhf0hhjK7CkWQaW7Z/WnViX36hxnoDBn1/3W52kzYL2VrBAXJvmkWp2RBeMi9SAfe1Tpb4ZE9178
DnTb9UUkMVhf5hn+k5H8baXUjj5qyniv7EjJXFyQYwc6U9Nchp99SdbgqgX/bYpNXTu36VkxOoCx
A+YsIBoMI9s5LbyN0G8ENlqdfkKlipkk5QCUvnUaMjUXhN9hUlA8SMNtXWB4y1Bh9HQ5+Wj5afxL
bOCnB56wdI0vPNE6OxZ/RtDzerKsTGelxrxvsHvraub/wuXwssnrtl88/zF97WzQHxymENfpGXtb
wDLJ9pD1vfn8BH0qap3cEWitzSB93u4xGRQQPNFLK6F7uSKZcRrfrzUGrp7sYsVMdbyxF8zMreV2
HS6v+41SYr9Bnhxjz5BbG61V1cW74SJKvVSGCJlXinc5DZLbYz4oB8IrN+p6++wlU0EAJVViS4MN
M5sSFzwRP1XXRMU7SSgR9tujiglEXKfcEniOkFHATmeCCGSW6y7KbtRL0L6QK8jRyB8DjwXN8YNM
yNQ/Em2JOcbgvVuVg5TVTdUfm3PmC5uPNWJPHMyT+kXPCUxC+QHRrzeWnYf3MXTKageYMsuIfEGc
+38XGOyUQ2H4unv5tpvTg9cLq5YOaGjK1NF2pwhWTtmtV0WZlvkZL+FZX5X0xHtxy74ebP4VaYGi
B+NLWyf1GDyqXWVS03/lRDhonFnqtqcoH5FG3CMGZ8W4UWRni6y+Hf3bgtsxB2WD1JSPqL/fHm+v
+WrqAR9lsAeZ1b8IxAJgd3f5uR+BHuAWFo7I/JJRq5qaU0Axvn+73HleQCPb3C33ZEvoBS4QMZRv
9Bdn+7zUr5QcUD9xeaH5ChqhgAj3M7/fX5PRMUpSFsbSjtEY7AHcsnFh23dtv72/DFwSmyDkgBRw
z2pevRfh4nH/hBtj4+LtNBUdeD5x/mtoV1G55zJb5lsIqhItDhyRl//+5kPU2aK7gRT/Hj/mwQYw
LngyAvvRh4K0TIYGIIRtqdTF/B4r3iFjdQhc1a1NUackPaE0G6nuurd+81VT7dKOmU4lE71dJBRr
rSMpmSV9tFVF0VcjOD5GR7qNw3VwGO7hB38k5v8T6luFlw8YwmeyV3/AUPV2OjRcN5ozIQUzCnYF
r6tCuWvjIcBcQDqJVnDYeXsLUzEkDtPwjayiJ91aLWArPKZTpqlDf2Gnh16QFjeP/2C7QvhfgB2N
LLpx45ry1dTt4o0Iud/Px3NlZyESezPOIBu+n1FQLJM2e9Sd6eFTbD+LvaH5d9t2Mkmq76a1WT1c
6tBME5FTkDvB+WfzBnDw0yAj9X9veLlNqkgtMUocMQh4JwFIPUCFNOrqfYDOaHSWVJrRovBKjZ3+
YN5ttf5v8BqCx08xwX/26mDEmFfGZE0KPX9nQ6tWTWSuEGokW4S9BHRos8z8M/8eN7+TaNunc4yb
hVUXMS6vIJ1sAtfmqErSvsJprn9Dm3c48VMUdYYkHb5LUI6dQb68TGrnzWWlTUvJWN4u0t9t4LB7
AcqD7ZNgtQGJw0HDoV/dAbG3abNxb8SDS/aqXUBgZE/WHxlX8DGG2LhqPcvhv00QA6WwvWjsWH1P
pISSy9ECNhGBAKnm/XBezy3Qg1GYygocgz7L3aPqmB+4xnuPsiYqIe8/CIHPTJCcqHbT8ZX4Qsbr
ngwmQzsJHctklxaRTzph6VoBWdsbldnOqGeAzic/28mJOvPp4U1Vd2VX5JOT9xtvg8RzdLCrsdYD
laDkyLgIAPhkEw/nhtPIvmTovX5KrH4jYUYnk6iRoh/TJ7ru8sB1WGn6WLXWcapRV6QHiEcN+dHE
sFTMEjeVE3iQrcy2dDr7qpLjQrZVRsh7PDZrTwgERwku1OrXCxQO+dn/kN6lTdoeVL+uleN3L0au
v8V3WMtv/2fPKbQYtU3Jt5r4wB/riyWfZH/x6i1zkpUDumsoO5Kii9ZTPSPxTx6KzOsauG8KaB8U
ONptW4T+8l35Heo5gUCeuDvQ+SF5hiZCwPVaz4c3YjP8BbUZcpsb4YziL2LzH2Of7v6t+8rAwSeI
DHZ4IMvt7RqgjTsQgFLsIbih2vT4n+8mpom50MDoU6JnWt29MlJFpaNcPQiFulGHsQwBmVNGB5QK
C1aeHdb/EbZ5jZoxXue9l9luGNFCYnvuKXU1nAGmqmsHRHvMR6S2J/oY5irzQgEBH+jJZT2YdOML
VxWHDr3o6wfXLdP7ifMfJDPlvTjsy+KcG24iLm87x8RJbVkFq+eNc9MCpI9JO2/5IfijThE9nzLF
U1L3u4fGjf5VQ/1+nT9hqGctVDHIYHZc2DPdXPqjZBJ6DtUzVXg6Qi5jl7wrH/dsIKfk3Aohmh+I
drBFzssV+tGVzXRwxyaA7i7YUkEH/Yt7S3OvkUDEvezXZJ0MGsFvQxBSKxkepA6lb9h5x29CAfPX
WNLiCPZNrfyXOBeNMu4lS8rM+8LOOvZ0feKShAILY6V9IXS7LbwqnIO8+hpQV4iTgAf495R9WYg1
7Fdh9sW4lzZ1QHgljaB9CFydlTZjUYRvfT96K5UsPphekuHW/tnOC2WSCJOBebBgG8II7yATaiiv
n1vjx07OSv2ERufqkqAr7KswCHS81DRDpRxbbUVazpkNRmE33sXOXJUAbTCMtUvDpGnSXtfTTjaR
5M3C66q4wrbyDObFQ8+ZjkYhpwCd9s6OKtVnwrFG1PIacmTZlAkzPxPt4ZY6oS6b0QzEP6rAgp6s
Au8Tldabk1z+m7gYEvCeW1moTnavN0MDz+cMcdcvcXOHBQGu6LG2VddI00xWTy55018m2Drz0/6j
Z5gjuxPO4sWB833z+PnkMFaG0krUiY+COyNRf8sox5xSjvy168LZcA5+Btjouzi8esrFFAiG/8hh
tQAVvrLM7CV76zfqh/h8VYqeRw0u/5y9C+xIZL+wwZreLl8OAlm0bsd5wShJSbLKAg9n3a7WuEd+
YoQvpR5xjha/g5Y8SXI1KjiFaOX2RcQaLNP6d79M4lC7x8o1+Wj7YtfZhJTpve1ZBpEFjeIlvzDY
bdJjsnoJwSjA8uwHgHdZo6QdlhiHaU/th/EA1VNMBISDISMLAuTJaZl+wCPoCh6b8yB657yTHfHm
UK5pOj1S/b+4tLvea0rBdsn8mCb9MIQ0V/cRcIUFaNAYAJmeqZD8wekKi9LMfuBnXP9oTmluDo/s
g8s80yBJEYi0RLBLdCmMAa1iLmqDKvDfF5a99FBNouptP65Xc2OUXRnvH76GN5jnhkBR37RE8wRw
DWXI2Jl45Lep/QWzqXmZwDkrS/uYOa8FltNRDy1NB+CmEZM9IQUN5V+OpmYqmV/jgeymSZJzqROp
LOaBJPKKzNB1ylBzPkf6arE4+M1zWr9WGcQT8qGCeomWkSL5rHbgmNDIPChI2XtBfLObFJ5JsK3D
861q1dqhy2AG0os6mGYw2hOSAsnjlXSrLoFCsb/KNTwJPVEhQH4WRNSviLbeLJxyTbQbKy05tsJy
pwHYG2bpE9nEpdZr8slHifvc9qvmQ/R3Z0PYt2VI06MXr36mXQApH/4ttlewYWcoXEn768Tv8ePk
rVU0gVpbe+Sqvfz6wqy9X8b22skYhh5ms3qud2M6KycoXiA4UMjp47aaw/NbN56vfGGQlazYNs/V
9b+/bzfVsw5Nhua4dQDSjwuicrI6rFi5RPnkVRC6Yu9cHz6QTqfDhPTaBS+Jqj/CjM5olrJ3AULK
DrRlrdzU1eaR7sIJg2RE1PUKVwif1tB51IW1s7VmZCppIvPAOg+NB4nObDVbZkZrAPaoPdmEDqEW
iG6tedlSphWd7Z3Vww5u1OoILs06t8fN1iG3Q7js89Xj+/1TxSdU5R5CK3K6vmJidfLiPXeHSnBd
xgM21k3EsagYkJBIkmk7d6UNyb6tuKxO8wpiQWSqKM/4b0HUNkJuXLe7PrhDPThSitboUU2kTEDY
u6vd5UW6ryXBHy4MG7CeMdPY3Qf0J3il2HLw3dTB6ItEnczuisx4KoWO5oCbFr8oGNtHA1TNxIiG
lQ2JI6qJN/q5tH1V5PgE+s3BlDirPAxftr6vkmBmpCfVFkS/fWfBKiyCgy1zxaA/xKvqB5S+QiGw
0zD2ps6KaMXXIp1TBITyx8qF7ZHBVbaJ8URmsIQK53rCQLUZAx/HsPrflQYdpIeGs2Tp9utC3+42
L802YBcB3lGFWdkeY8IdKlPv6YsZxSmcEQ2R/WcGPVPumNXpPTlqQG/o6amITIFnROpYmjMPeC8W
/EUwZmm32X+oXCNphwKvnt+dK47YnnqdLpw7eMzIbGp0jZzJOA8d3XA/+leiSAGInJk26Hxf9do/
jl6WBiVdqwoqglWlCho9Ik7KM/Wy/GHsJouWa277xP3AHstfgZNwvA4nISGBbtPj5fsO+v0rawFI
QJeCso1sb7ufjq6hFx59lkTUaHDIXVRwTtTalo03hseVWu4IOfhmsAzbmD16zBcXDSxE8CtB0XsH
XQXxMt9OYPm37XjDoHCT+ixPCLd2NqRsDXi5y7VmXWFY9H3Uy94pvlMFMvLBIDK3imxaQVUUIFf4
7+XZuCDThN1y00ygWAiFwB81AL61oR/KQM5GOnQG2+GbiyJcugCmdQ06z6x9SSKMGLVQmDvSPUXq
EpYhWzuNrFIqeew6X2QD3SCqSt+75eSv1LrnltouwCE2X1Z0aPfPJ8LkYUHqLRTwbq5ENYvx6GRk
Cyd5NbMbbIpYiHqO3eaLmdrnj5jXpcdPw84BKUBzA5TDcE7I9S0tzKAXwoV6JDMYmk/Smf3WuU66
DRDUA7prqDqKUGU7ABbV5UN6zjGy/6E4J9Pxp05uhbXaChHgCnOvZHJ1o6DdUJsPPLnBxdtRbt7O
pXK4D7uE5kA2FjM1SKfuamM++lCFKQgN/ODdH6pvyvgCRXaRzJONI5AjHkuTRPDRTzJXHMLNIL4f
L/ZR53Nsi04NspoxudBxr2Z5LdNJLUD0u0qYk2Vxboadao6XaBfKrwu75CTcgE0NsR0g/WaCkcAM
7YtatPvfetCZfehjbmwm8ft/tJulIc7BhMvemlCeb7PWJyaoaaoxntC9Xnrm2Lb7QmhWQoDNYqE0
faOzJgwkI3pvCDWu+rcxtEFIs5IFQ9mHTgQsEdz3tTi2M27eIWgrXKndNPjYNcHL22IZjTfjjCcg
eGzZ5x6jDD2GD8H2tEnmNj2h0L3ivT68Zw8BIcJhdRGR46+Xyi66oRqsKySfhXcSZub6XdxebQD/
v1DULULcs/rQx/VLAaZw4ThNb4KXlCZR1hBvKmar3bZ4m1JKMdXRxxZoHVAK6NldTIBNeoScp9yL
QqUaeb/58Lm7jCmEbcML6DlfFnrgSwcdiBz2KafKW0VizOxVn1sWuVvRb3KfVUFG0du1eyNlCCKE
SBzvAgnxfLRrsgjdRPlzm1EqiO6Sy+hJMD0ZQI4z1dDxmy1jctsSBkLZtnAlebRaylCSPMhP2VXD
zcAGwzEX+nXuUf5TSXeQK+EGDBa42KrvNdesnLtnH/VGZqEGDSouBaTEsTldJHWplC1fI+P1nrkX
v8H+W/8pvebWM97ZMh36vYJr5AyjO9cfmFxZs0pbgJWCMtwtdFhwVVuDoGRfhY68JBWYfe6rFOq5
6vBDa696Jb3gnQvWjWoQsokvGTO8Nh3vS4yg1iIB19IzzGQXRRXvus3X8tg4ElhRuA4ttSo3QTJz
dlhYDcAxyujHOTC5nZtdVBDrL5Thex+FTRq58nKR+Hgig8d80Fujd3MhtVqki7FaLraN0KgFM3fa
P8da7xJ5dDGA2A0vBDwekzf2yt0/OL0Ie+W6WaaesKy8YUQt4/+hRDrCmfFy1G8mcU/8i8kKumMo
5nqlME2aDV4Icl+Lz4yBR7ycimQk+l1KQtxzIECe0O36VnmhW6qlU9HHDuawla6jctFim2Tff4Ce
sVwVT8XbjUY6hPUWV87fLlsDMhpP1LGo3/64EWSh/2uMcB5MkReLyv+OO34P4bjLp0VhlNzS/WBi
YiPXxBq3S2lUSArILSHjPzBvlhAUIDGcONULmh5nz+Kp9Wx61Y6Ck49382crXjuW52ezuj1qKyXN
4QNdXeyUccL7xXA7ttAK95bF/jnMvI1VTdrYgs701eUcdBoS6MV/JoBdA0xknSMNNnTnp+2JxpX2
cwrr3zX9zZowRB2mtF7+UhDOYloz/6ou1E5OBTu2fNm1HaZwpSgf172VOqSCWlEc64Wm9xBoQqp9
RJsdVwgF+nCnK7L7gCn/tLIaJy3smsm+n73UqxYENu/kv0rd0eRzRMa5bJlp6Zma4v8NKqc+Ynj1
i0CSbavVIKAbfBUiaal4SLrw1jIyvy55LoXjSzUGM+YWsvgFfaFOQRTmUX1UtJWD0o+eNJ4t+hET
+RmpPchuQxPo+P1wQBdid50jbdiU3C+ipn3iB9PsBdEteVXsmJ9IBGQ/HsrLRcnIMNRY/018+SlI
WXmpDMVhXojdtWNfAFnpkfPDqvEazLLJe5XGivyOxKn0SGyr4SKsDAGtZzghLMkPR00I3FInDgBj
peMFSqpLbpjTThXnzH7CFJAURdTklGj3FFa7MzeSloZLRPGQMc3u8ShnkqC5X3jd1652EmVF6KEk
h1E5qHGeVVP9PxFz3nnetj88Q9Lu5DpqHsFt5qC++pG55uuq9jhwuJEM27XvhgK8roxewCrwGJtP
fxOaxw4fuqG5/aykFT4+yebiGpkLIA3Cr32XZQR7dWs6fFfujyME+NEMTRQ3NuKpfAUdH5Q/jE9M
MS9KMr1+NFPqRyQMRy39vwcwwF/ahXauWjP80wUNFr0PMWga9IxpnTNjGA5b8fYMUSAems1vXQhf
qUsuvZL3RcSUrAILETmBRFtzEdc4l1c0YQ4LHgJ1nXPCEvlqfTgoY3G8p7ZriVzZ6X6M+NRXnMhw
kDxMEJ6HjojhPj8ceVHPInGKVlY1GjkPRIcVrpH8vA7oQHrlA19lNlCQyjAkXYN1GaTDwe2q79Xg
8hX3X5Pf7kLzJwPZ/A7TUw4LaaRXe+GZE8YaMuHKY2cJfYZGamNO4x/V2pHR4sXx1/gzj2yYK5Oc
KPca+oFa8xfvw7vUU7WSTdbKJ5L/Qwxb2PHo/ysfKPcvYxK01ASJNgSFf7o8Kswih3QjRyCRNsUm
3NiS7ywe9APglGFaW/9qDE8Nm5MBfLrz8LNHVvCltkaWrmH+WtOant0w3kl6q5RDktaf4WUiI6pS
1XssykM3zikwBcxQxfJKnUVLednxondmt+0RtsKOE7r3I5A/gmpdlTHQtXoh4EknWqiADuk5C9a2
h8EIGaF/p7wvLSIzAT9aJtQ3QxgrZS3Cm5qGieL8Z3lhTjwdeaHvvZh0WrUBLmeyjYkZqtd72H2g
+rOk/XKc3QdKdYfMxVIpDiorahjJaAANbPSjXERSmbXWQwwXCv3b3MgbDVeiZyw/zDap84oFbiiH
hhtPu/wOCr48Y+SKxIGTBkFkzIl84ddsjC42GnCOxeD/CiqvTkYeW+DaqgVMSeulZkj5BTdfimvr
coGUTFr+irlTUtnyBA3rxaVPqB/qY26UHNt/z2+ytJZhYoLKnDLLbx4HRRTdoQelIFJh62vQJK6K
EY8XtuvGLY8HH6omxX+ZbsgM9knfotFU4feb3nFp08fiWMelQCZH230qotmC7MUO2WXiwyEX/1ww
wnFLiCo6Mu/ZNwsXSgoEiRjcpD+IvnJD5Yf/0e27JckOquo3QTwTnjnmx09UUG6Q9xfyLe7KzjPM
kIL3Mi/jvgfFRMJ3l5aAv4QwMAeosWB+SHn9XpJinASaqoE5vhbx4lmd/OUfm7y7tDJrC6R+S6NY
KajfUtGp8o66oRudwSQ5MiLSlJoUF3LRVuPI9CRq8r532C6kjlh7aIk08mIl2V86QxubjuTJGJv4
MI1N+8JSTv5nzh1qcyIN2r9yh1VJevWwRoeDWEJ5DnBV2bnsZskB/sB/kQRH08eg+xds5SYk/c3X
WxmccUeLPpNtT11mx/GldWMIeABSDYoegfNzPVoR2u/WL3QWjc+cDEFX/S9Ml96HHzUApG98gvnT
fPybFweWcOIbsN7QbZb0dU6+QcT8L4/EPOAGZT8xZK5HzTgiLdHc0FmkjCnEcUzVV9yXr0CIXgAS
ls4Fv8qaQcIsDsAcS0SzKJ5gwO09IXUEmFAwkNUy5giyxms1WVQQUh4L7TC3RyzBcbLl915OX6h1
fXY66cx/xhF+R18sy6QQvihihSHMtXRnz7/WKPjJncw5OtdRav3vImxRT+CXuFLEyFG/ce12jdvm
gTBI7O/bIowx0GOA0vrhdW5NOpGgzheWKuPnoCEQuyMsb7CJJlwAZY/UlPrrp1/FsBsg2q6l96Ei
45kClrvS32Q0ucuobauEZcRY/PHkZtepZW0pV9RBiyubbjbfFOkYI6176K3ttJTlt++xrlg5nXl5
NsaKKYwSg4NVvgKvErPivYr4pUezigcJBL4/ARfJRU0znlNE3UAw59rMJXHrgaealpcKXU7bX1DO
UenGTec7cwKEhfK6hYegINHmKo/6TQ7JcFeualk2hxeXGQkYOX4Co4r+xzFU7ae+DpZlpzRf+SCZ
iRSOIY40UHBooxR0J8byn0U8wygyzMrkTaeOdbuPyT3KqCtK2Ctyw3yEDmG26IzES1KkyS+xAp7X
BMwzFj3TdO+PuFJ6vs+x8htE+FJTBYMIOMZnue+XH5R2y6OIxjOg2zdDs/SVg7DGzsCQenJYpyVJ
kEz/dq3p+fbG84QwfAxbZj9P3ipNpwrKeQULFcLGKMvIezrCdM4Z0ry0UV2GEyYjJDDs7HGXCO04
RAhPzXcnTmbNlQBwf9b4hoVi81lw3UiauLYLLb/cYWTLvZbPVbZZSLKTiR6szNvMIJyi+Bg5oSra
LE4vQBNkshN1YzzFobSOB1CBEQ5ZbMjfh9t8EHc6YsB1+6X0C7m5nWamZ+rxQm2qZskaCjH4KHvR
r0vvNsMjLPXJ6eFYIeaVgPp12/YVIT/827y6HoOuRDn0o+t0hVouoWSdTKODxSxsL9LDyIuKs799
rURtwt0uQE6hU27aOwwlEgPvm+jA3+6mdrW7SFv88e5LoXBr8UJqa+tMWeKgmWT/9Gm9PMviNvZy
uW02ILBd+PHprpXg+IEClteGrV2D0+6s+p/Jd511cHl/Kzz3i0X71ekq3Ovg+E5txz8InlIYonUG
G267g7LgXbgyWI6rhOBL4ub/o0db3dXKAZFHJrKJndt8szQFtcUOKvYQq0G6I0arty8vmQs+MIg+
2c0HOrAWWpyaqb67dBprCq1EKS1NrNhNNln9uhSvtDB+gtIHImManSrNjpIbJnyQBPKp8cW10H5b
yWqxsu6kl88b0aabSSXK6y9edtDEGKnz52nit1a/WI1iOeeSFUJ75yDdAwpfvpVflBHYYbHrpnBy
RkLkqpWBaYOBun1fm9h7jqItuYJrBEaZHS2a41+IUXEdbJYsl7Mk+dxjSTJF0cOOnpb/2uyotAlp
CGgr7GxcrBZkI/IUwxpTgvRCySp5wp9sUJ4NVcS5a+pw7e+Ilsr17YYHgUXhkJdBYTnNI7EXSnSZ
+tzhOt0cx4RToE4GJvOCy+//6vgVr1BCZ/JZ8T1GcoPZ/16BkP83sI38ceI7o3c3p8IaeufbTJqI
ymj4QHbpF4Z4vIVAxxEQHm3spYbG0IjL6j5t5okkd9Qhj4L/lAPBniDwbvrc8WSNSGU4rZpxYPjc
oZMqMfEx9uMI/7jsnoQiS4DSJJX8VymuTwmErZMpxxu86abPrq5bEYNh/8qk8RXe+akk3027j7zK
2sKBac+VHZXVP1enuzxl8t7wApoGQJ3eSOnpXzwYdpvr4mQQjYOrWN0NQFWdFqHrXqPluTv/bazX
idQD1wSqV/WBTQATNPJ/4EXBHIPm4JNaZQ+WdjOMV6QJbkq9wlkJwADihu2pX4dDOyEl73w0HNy6
0+xh2UPFPR2FmNaxpHcKDoakRmPkhJJfxyUM7hQr1mn0o1YYmgkodE7zPRQYlbiKWjwZF95JA69g
w/cvt8QBaa+eGidTk2Ec3qSeK1Il+VYdQx/o1qebVztufyDpjLEbr+rOJK8+Wwx+HCtOFTrkYXX4
ZZpZk+xOKe9AWRuOIGHZTQzltwniw7b97LM7QFsJB5eOpA2MIw3q0QdxLqlDWbUq0zwfaK8fSBuf
YqWocxeuj1G2ApsBZF+tCoh4I+RvMF0STnLj9SpnZ0NEU8sO7kuJ979G1vhH+DBzH/7wYzy3VFVc
CBMqNtF/wWTIVvmxhqp0SNn7uma6otg46jsOn4z8SEJTEeDI2JngU3YkEpKhEgju3br9CAxuWi88
xJ+1RWSOEOfwhXVfDfS8tsDqka4b9NZHqxLHLUEKDai+v+PKfhbKOFU2bdVp6twpPOJ3udF/2Tn9
AEZm/VNA9vltKYSyDdZq9m3Wz1zHIO573I3ltle4kb0xCCF2k64+oDtjT14k1ZnfOIjF99DTGXYe
pNrw+kOeiyWZmubcCjfDk4XsSu8w8dPVL2e/zXAiQSoz0nJGGWfQuCGj/NxhIUR4w5ujtl0q+pTA
PuTHz2aMgj97vAAkDX401GYUdhMtQ3BVFDMEOm/bvXbqFGJfweKlvLJjAD4doC9OQEFbkYb/FPW9
6BNExFkRrQFuqNB/HUH61nAW+ehWmtQpv8j36xVLS2Lr5keuTxjTMvkNAGop6AQlJ8Ent13HaOSh
55EwJTXCpXdWACakKabX17EI/67+k+ZTFF6TwnygNYFemeJnbW5qz6RAUad0yQPhNg1dVEx8lMLv
5iqCse0c3zJefSTZxPvI87xCwHN+MT/eA7SWEtDlWxCvga4fTQdhucErr17fgdJiFkPa6aLfX/ss
Q+ySWKboQVq2jrv0k8pz3Z9J5oE6sKerUDipSgUddoP8B1hmtvU6PYSl1aRhdCdSU2EWuSF5954w
ysXuWVdeTgJOGkLVchN9Jao6TIjwWLmePdihUzTxYELAD+w7sy/Of2Dkxix8Q72KcqleRKbr2W5N
MW/JhfPd/vrXd5uU8oU3cQNq5s/yy9GAm/8VWJkv8/5R+q/KFON5S3yAS9XmuVCJpMwXhW8LWIi1
hJeAUW51dFZ5QNzdPvpNu6Hcb9kZbWXEzSHdXvjBXz9I28MdgCbRSyZTWJ0G6CR0GKwYlQLznwJJ
PtEGOnIfTQWHGNaWj7j3QFckMRrvPEHgOvPm3JckvCUW/k483POso2sISqpt8PW96D0fwiu71Qdw
sWAPTjCW1gwdIx2GDXmhiLSQ/DUeO1FiLTF6uH8x9364ps4RBITI3d5EzyriNiednMFAhs62qTYD
+GIdxz1M5pULXZZ22BE0TOS6E54bdmTUD0UvSx4pkAxs/2Atx4kpAx6DcnHLcuKpDpPQR/m+qVya
b1soMUhjTX04s2Sw8jKFU3k6xGfsyQ2vJWX3DtEnvfi9yKh+SFUNEU6JNkdAmDZrBSwLQ0ACII+m
tdWugLSh1k4lodFveS1G+55U5SakA9/HwI7eE6eNwRkLbXlA7yRM+y6KQtDwVnHoQZTEuofHtUbd
UtKzb566OrKsC3h8svPmskHqfw3fhjqKw962Ojxd3MzwxG7vn77erbl65DOEB8Ac1iwmeMANkK+e
b9xhtu8yVIneGR4uaKcGRQHOjvn7hgR045pehq96Z1PgyfSuPYjXR9ug0WpgLyjEGxeH0R9Rwzp9
lt8x5G8ecuHXY/tf5ttCX0h61q96xHO83xKMSQnEuP57Jwp6cgEALcyLJNRDiuPa428zbw99z3G0
dTSbYB/vqODy5Bu9PlHOpHwCTUcWhgz5GuW4xzR5trUIe8PtpuN02qAF5eTN2c/OnxEOY6GiewHR
uWBsb3Wc0QRXGs4mjUBv27lq0msBhBMhj1b9h0MWfUiVsCgpwLWiV+jcSz6KWScze5lLUFyhrz/n
YAZLAaJbjcE6yB4weS2A8eLQVQuUV1GrzexQXIbtnedXvoUAVex4ZiOygXxyxjZR6PzYoZ017pa8
++5kHUgwEjonr2s59WvCC2Xdc0Phne4/bT6pCfT3sbPMpnnnyVyZ8rQa7wggRInSpkuEY9uITbBl
almMaQ4IPaPjR81UvscgZyZb7Ilu9SIkl2eQtWY5aogkwhQCBspBq9VeVapJEjBcR1YYBmeXA66r
48ssA+rfJCtMrFsmkQqLV5QK4hcBadkiRNt65DhnrbzcAENPeACpml3lfw/JgAK8OSW2BQ8J24M2
olVR1No0NxoKyuUiD95Xyb8XwJD6evAfYLvNA0lPNe9c+pJi+qNTXzgbgTbezskz76weLElzLzqy
d9iqqWBjbZ/Ua4j2D7mj0mhWhqyF/w3dlNKyPWwHd+KWanGFR1gFKMxh1/+NdEK/OZnFjMu2UcFl
NyBZJvNEgQCB1/SubJM/qS9r8gEeQ3UerW37gon/rPYUSAJFbdp5bp9U2OZzH2X6FzOQGFvEL7T4
UUXoOkPCRuMOxZz5o07HiTK5XfytfSNGT8pXy5BWzY2Ag8B99MjULnyMltmG9MJwb7AlCyt3407c
/+HmVUbpKWMRvoqSqg0NFNwjAAifdxUhoPA6Rz6qhi+IL7z2Ksub2hxIDPK2Wi8LgxP0nYonitnU
M91OKXHRNAvthfIidKO6QpDe+qTDE6WqduLX2h0+Cqwteh6NtBbuiGo1Udc+eVOJXaGXRUSXZJXj
QVhYdZuSQ5O4kSXZh8uQu5w+9J9CHrldOomxm9Ni2HEIFDAfP3skeGtXKfo7dk6+6ZNg6hGy3fG9
Mt7cRlsDEddhxyhr+t9kmidbk11V0QWpe72bwngyeCXGTHXh2ucg05J6r0+QLQY2xOxoVx31agy2
X3uQxMW/UqtqswF0PyHWmHTCyJM+KfCtJLiHypWaazgRAddWzF+MxLBPjLW5f09w/7anDe5TTIY2
JR/uN3vyKW3PLiX4lopHMUPN1sedW3Ez6zQkwQapvdPTx0JK5q/INtCBVrIfse1Ifr99ubvPqg1F
ug/8ewilQOnDgv7JpgkFGGGFy6KA9pp/6t3S1YZvDLtwJ1to9LVCS1bpHs24p4ASOmupEfGpPjs8
LzGwCB7lUgyke0MWW8F5Z5A1SaZHhCdro3CAqLBLRyif5QSWfgOkABX2sAxEsds5ZWnZxqyWvJR4
dX57ZcdIi3YLa6AShCGXSg4ErNQAK08PTiibeFazs6hiut3DiLuJ3a/1N24fyVsQEyPu7PIMxX+p
vWUliO7hjevIlSpIGD4ePrCmifrf5f264aJQ+EmuX4kNR+aHq5opFY1ooQwJmx4BYhzVU0eugQLr
QqtwCBDGPxrf1r7xI2vwrb5EYxn9EV2iXafDOIyT/Cm4RP/cbD1eiqdw1KgUvh0PxchJu8XWX5Bv
CR9G+CGhVe5WsL+ic3OpdsYk3aT12bIdUcl5PY78uXMk1ty74pdvm3fV0S2/+BHGqqbmQ7L6GDDr
NsyfRyGscI0b3x/CC07Iw1QbDReE9kPaCQGFjFNxxaeLK6M6Qj7sm1N6o9mVirlK0AlYGGdfByxI
leWclm7JDU4HiLXCUle/Qn+hH5jUD7e7Ad8/zSSiT2hEFO4vnJ2wghAsP91qErR/Gpbp5cegDHks
7e+U/gwSe3IcdRx9NF7Lfi722P8qd1VqJVC0d62nWisZBL/+seEEGDV+ePBfwxsqW+Cqu45K+tlP
xr9uyCspKelgprqu5ra5SJdFXCaSvp9HrphI4ImIrMfBdfcy1dUHKvOnGLarYY9G4E7t2LzZ377K
j1+lJxtmZhs3btibqwTIspcQ0JBQ7NHNs/z2PWQzfWIYnMDRMabZNmNC3jVNqGgu5oS/hiH/PJMc
XT+1KxmdGMmz23HAb1yRPy7ONHseiJkHYKXjaiZEfS7rpfawZ0tqISmCcb+oF36wcteuU/IyCxoH
MjxN8GSIeE03CpW34gN1XXyx+eAKz4AqruwF7SFrAi3lRpMYBLstZodYxzpKtBnzsjZFZpHqvpM9
BMqsnLYpfDvKDEMLWHWog5CyWCsWd9e/GD5LSgXW8eBUhjhFjmEwjZEdeYkSWiGj6ULmENH2cUGK
GkjR0eNaJIYL6FeBOW2kleW7tPcpfFQYf8KBZLTvHQuGrVUZbyrahwNAx5dqRGlFaGD901h89GYU
gC7g3gowoeP3RIU5LCa4exQYgzwp/fRET24eRcWjeaSK0FojpcXEn2KFrzSFezN6PZQoxPmvY2D2
CNZS8cH40CPpCenjJaha3oBqV46JqMQzIe+A4KPyC1cxr+MsyOajHRiS1+T9vXRCXUKB9YUd/4iD
B++pvdfMmIs8OM2mQ/JN3OxyZIn9mhUcFpqcj0OXH+RXjEBy6xqClKIR0zny5zZZ9zxztei6P0ez
Y55QJM63504w3zvpaKwURLcKD48Tyz9TCQJRZ6cpyD93lX6IEYZ2pObAfqpKIf/cTdi2TO56g2xh
9sydVHSRiLqvKS8ADYW7MZwWcK+L7AXNp7s6DCMZcK/Fp5Zx62/pmClc6S5IG/4urGXRxoMHmrDH
VZjmimr7aQnWbbR8DXdjW4QRvDwhm2CXV5fb7pgu/+F4KOBdibi9+jre6QZLdjhIv7gbBDqQQInk
w6b5NZofqfd5+jXhwOMosGUnMriX2/plXWWyCk7AOobOUwm010/NK1CuIE2v+uqgh9poGtqFeo7Q
BGPO7Y4kn0E56m6iVZ/W1caEM3JmzOZW43a51/S5fsn18VsZ6Ld9/E5bNs/CjVtzTPvdOJgupMOJ
QV/yfvMaQYJl5ouhe0OV8R+4SgD6NPg5YvaJ8YEhAcEiQ6/qxX0XVnnK/JSGfn+qFmiBZQU0GthY
52F/g+XnNlRGxkKwxao5iKFAJ1qFTgfFe3ytciBEYlz8HOPMr2ikxfLYOJ9+cpczfjg/k1Jt70th
F6U45jbTgfWzlUbHcQt5n5ZSZZboDCj+zvxKcyydxMc/PsCHOmVdV9L6OEEXG+u4RhX7gzQfgaEy
wZTD2uLLXiZIeFaHHJdPfpMJypND7NWuoE1sma+WWXjbBIgIRrvk1ivtjgJMA74VBIyatfolmIus
19bFxqo1YpyTTZCpGWQKRY1GJE49BlZnxy/noX/wC6s7sJDmMz97dyXxM7KNu5Jo/tMYvaksqHuH
u2rnFPUXENuMQYyPCpGJxdeGhvOYyjs/brK+9L/IiRaV7QlypN9AGXPPOLLPsJEPMksRYYlw3AdB
s0/5UGjs+7oOz9sqiH+mmFdZSuF5/5V5cOHhTmtRn+RNkiGXmz4yq9iVOFrZC5jaAyckdLCJO9ya
/P5COhlF83TOutdsTgnL+HwFFQA+aqELYAiBdhiwWhaqBjfgfeacD/1ZcT17MFIY4Ecr9Pi9Eqt7
N8osZQ6jPCedEWuwGYp0OVu0NfWz8QYFDyLA/weIOZL4gUwN9QqEuHKVsLRdDGhIkVO3HEbSjYz3
5JArg5u6MX3VV2b97zRAWMSKtyCVA/16pgWV3NHGkLMX3mvOMBB1aEGbMIbX1ND8/Q7ZOjlvU+5L
K31+oEkPEJ5h8mEbIvT/RXa5rGh1bTp8iu+uu78uAFOZELoYxQpd6vwmZmfP6Ze1/kOUMIb87U1G
GmfDPJWDlcVFGdFlk1ZhLQn+3EwNgQAi1eVQZlYtjHcE1Dqh+64fW03G3zfZkUL+7xDLpOdw2mjb
7+cxC3O6lZKZZPFI3gtArFZLmMGHwx8w1z4H/fLbYQtEKSLy162FHGbPBoszbAnJr3k5OOn2MVYb
pOZk0BsDuE8DqSr8GFQqyJXSAX2H0ZHP6R7sbJQQHckBON7n87tZoIUy3maSYQ8Thjg/NJRppBda
dPWwt4j3qhQZeLUrVFvpg5opxq3m+FHNFftq4qVuSOXNC5lBGjCnyV+2gEcQdPlaCAADfarfQU+O
EQiCjoNGwzX6+IPjfP2/4EKhhPed9GtZyyqkcQl5sMf78vocz7nF4AK3HM/o6eYmpScojsdJUfK2
Ns1eyD/tmzo+4CUqRsZajoGPRL3rf7kLUTDQ8OD4isTzwYmbHrjiB+op8HRKjDd3cE81Bj+hQzBR
Icc/Av/qbNpDiCLi8KidmBjp+GYRFXCO5bOGgbIGynODNHv8tmYsLyJYOyErFvMhQQhtcQMk3iBs
KP1cCeiX9DS2W5vqc+oa/FaWdFLnXRe+jw/9jKM/Vxb+KnMdsCWKPe2xLoUzHsAKSsgNnJrQXPz4
PvHyQ0VArgh7a6WOMN372qQZLiOyV/aUoCR+SItOuiG+OMgfEY6dd8gE1b0umH4yDU5BBd/7Z1ne
A06Kwsp+GMCYRo4Gb5OVbPo7+/hQ5gLAQKPYA6FbvklG76JU9l9xXqE+cLpdM6ZeBj5lma4a7Bpg
LqFtUBkMUjD8K38IFjy1KLSJ59oWVOYSKyEe6bOeWQudi2CiHmtbpfWWRzLAiMwI9oi81YvILXGg
BS0b9UGrOt0cBEA1V9k+DicsYg8fbULMiariQgPP4GBvPxizSxZEiGn/3M1ehOTkeIxxT1egyHw6
dT4gbSRG3uf7/BguvslK0KnDPqGHwZpEd9RY4S2l23TY+t01W4k9iRYXQRfDlQ2jWgmqhUjhsW2t
nK58UtQdNmcHH/iXcc0tCAyBd4RXpnETYfnGk+v8C2eaWB/tGXwpVZK2D33TFaCCw0JtaRpoVhCb
BQVoV+lpbfe0rb0yKr2Kw0v+AydDW8c6yZf4H3/htdq5biGFuayk1f8aaO62OEiin+wwths+S/oh
jjY4j+QrNasiF4DkAjjD7aXNCaBH+FRRRZP7Y76VJb5c7z4rq96AiRatRwu6UNL/QL7Yfbw9WT38
RDY6gTsoqXl1LXZqDKJkAFoq4QRXon7pmXtcP+qwFl15eTq1i3Wzh8pjrWr8usdjVnZqkDtXapon
RnK5H7McmJnUMcs04CI7pDlfUg8M3n1FMKSVOSS6GUQTbc2GDnW+1mFICULSdw4JtE0+kNLeAQrY
F7rqtg4WXM8v5EGMudwnx81Y091U/6lH/8Bx/AVEjtcvBamZ198/R+s1Oj58tzcdyrrkiX3R61ub
KJeS3wyUjfE18WYiRG4IBBbBqa0c6+YEtbEDe5I/S26GDEi99fbJiOykBj07oFIUPa6SqnQIHBj5
7hnusTvAcZyELDi0EvEY4bvmLZXhigM6PFq/lJt2CA0jlsfJtgOdPrQfpN9xNX4KKZoFI5aAoIx5
qgow4F1785qGQorGAGGzcPjPCkPTstdF4i5FZ9ybTo/NsIk5t9MPB2Tncjpq0Ur3NFEkR0Cbn3yZ
W4Gb5da2t4VgV7XrWJ4/mHgxr9a8RhM3NwHs++Pf+qojBjhmx+fVllvigzNh0+qoE1JnUUjw/Spi
8tgWzTW2NNY46UElqHB6xWyru8BgHT/YlkvKSYAv4YPOC8QA43s+N7EPYpypw7kPtFhVRt4NmvC5
zZQehgN0+U4rVcsQDmTQPzqGGlM94wAiRKPBYEcEpzOzE17UNpLzS67vlihAyLrW4X7cqAG0uJzH
7SgopdilWGTu8qrkbd1ee/f6BjrNF5TQ1YsZ+gqu4LCDgvWQBW1YN6bsRz2j/V6uKqaxM+ItD59f
7X06590iJwBG2Fq28lfM9ek9AGoyOh3BJmPHv/Nt288K3HW9rZ7xuIaBwOmnPOlWM1WAJFd92not
u5wRwiNS/EFxrrak/GEfn/3aPYda6de8ZsYwfatGjuDnKiWRKOi2etDvuiRcrZv8bQdybIoq9LVC
lrTtunZIxyXwDetsqAhK0biVBs8sjqUtqKHNSerTBy1kaP7HvUGd8utL6tbfWCUfcMyyakS56XgF
HPjDpNZYGBJO9DV1CxNPcAz8d9lJljOtwPn2kjwrFl878LYoZNxMH42TL48JqrwPjyVvlLILJ7HO
eFWqxyR/M55uVlHYKjFR8MkGX0811/AQdJZpbDjey2Zunn4cDMlGxKBJAW9H07lNZ6zHa411duT0
MsnMcS+l2l+tDplrC8pjbSsA1j/nap8KBxGkctj1rT9ka3eocunTGg1L6tN6ho0YSD9MryB1XyIi
UeivykwDMtB5RqmjMuPlc8AL5RfGWi+HE/tjaoMzJRfhxVWPbaagUY53mzYFm+NX+UWqFzR0rNmR
wkwQzR/XTdZLzxVfIVRgYhdOnwMPuLRASQV/Jgr0Ko55RxNOzyf5+o5NV6HGRnfx7ofioB3r2HYB
UbnhLMm3SIQfjB/klUk/urlSaymxKW5R7zGZWa5iTbey1VQX+WuK9x2vJK0yvCOoRopEF2CNjfzK
xcuZjZwJ9qBYjeHfFPZXYzpqdSVIRgjuC927/vtu/Z8Dt7WJvRGwkzK7dUfp5t1VZkqv4eP6JJvv
r+C2sV50XEM8w+LHR7QOD3wEzOZl9l3EZ5fnhZaIK1W2/EeRajYYv8vCcTuFVx6wbLaweGEZTegy
rBy6k1M9ltj/QRajK1kpij1eDfeEKCOf2oA7JE04Y80WRQiFOH2F0aseESyJGXh/jFi4+BIw6Hk9
fixqKpSuLZFG+CsmZ1vqkenVtBv5eJOxB4R6C4H1wLDCE/m4apoBDuEC1Gc9gsoPXe6x+yhlLoyk
SOetCyEkipxVE2lw4OJhbo6/I74+pSSP2E1UwTJ4evF7N1WFXtF+mlbutmb9YjCcEAnrLFQrNut9
ZeF5D2xOrLuhMlMMT8MdC7HgNS9tKB7UDO5ITgyJ9YGgtQYMkmTOYiKJp17q3DOHNRxEuUnjvCkr
PtwA6t0OTZsTWW+ZTUMrMnqDqkVh2TW6f7F+A0RLWHmxLF65FvvWoOIjXvgSvuYpBvXpP0+J42Wf
meyJ0NznH2kdFK0K8Qin4qmheXBEXg8HiK+0v5ue4tEpg1p/6C8AsrkNPztD+E0v0hztFCeY/LD7
0x/Y1tGZoZryab4w+87Qk+K5GXTOZOLAx6DqZDI8UKPMnk7zDOxEuNls9g6a2GGcJzGTGe+PGIpU
l1qHWzQt8NHrdbBtvSP/iNId/rmPnHfxG+9M7FAGS8mUNqj6inUR9I7DTW+Emcg9ptgmB9Dfej8s
rBLhrVJjdc1wOk4YiTqVgRtpCOWx7MJwDz3jpqhP+AI3xxmcQ0fP/AApkILgJt1rFIEUaOpYgHwt
mEY+oqMNrU+XHTS0+q1qTbKnoot8y7pqDq/2OPCTIOP9O6RWqvABp2PN0EfqVyRTcFnEOKccK6eJ
T385KLZaNFy99xHDmibM3WF+NeB78ltMJcUPIR8vnsMTGfnxjlaDWoBhVUVBf4LsIUsCadc6/hR+
6qzNb3LCvM8nwey+aQY6d9QpKbvO6qYMEKNGE65wrGzDwt88RVdwb3RG19JDwxUtHBLuAxnnaHNp
vacmH61S1VsktgmH/7TCj8tCpTvDOd/fpuUNndYO3MVBQ08qlQZkZyx3lRRJHXewALlqKgnrnHuo
mPcHkhRA6zt5FcykoHsI46/+l4DLQxilgP7biBy0IcuGqojpwUujdhvcgibv4jJtTiwfGJjSoOiu
4fpMQYJFUd46uP5wSIQ68/JNec6ecfi7CX0N6vTiWdu+1/eD0qsLz+UtL5wEgcxowFS5z/VYbFX5
gyktp4NXNePOia/lFEmY2CbN9ikXLRRsiN1xhVPojcheh27b7yDl9DyzFLvzjatkruHB8bRO+CX3
M66fA3gNpJnvI9EFH+0xipd9Tlesamyv0EMBV/cVKgvXEEqsCv2cxjDQuaGopEbp8XIFZOZKtnx0
+QxF1xEsqX5FDTad/E33fUdZSwWhVfeNqEds80nmPeVeMH6l45PUMXpWq66T8DZ62FZf/gKQhmWt
PbdUjNudUA2Lk/6eukH0zP2wla+jzq7sHHiI5+j3kuxwx2YRsGkqgSMjgSYIEVMqeUBJe1BAUwFF
k9IRAbrCyY7z4S0tCvrfOV0V/kdbyDf3MdKA+5SiVyM/V56MDr2gsb4WOXn42yYYVVLhXchgWVso
apScUuY4yrZ9mlf8y8cgStml7bi5+zXxf/3Dh3GolQZ3jX+OGmnqPU0b2l9U+7ke9SkgSRby6o+Z
aIIEQdkol1IodAX6bPE3sLb7M9Ke2XGi5UNi3z1Vd83x4tFbAWR8yByQBfqaDJYjfsOhhx23TwsS
zZ8dxvo9z9NOCF6Km8Sda45y+pcf7XyCL3idqqzbt8DCgEV8y4BHvSKAyigKEyq9yQSunzCQOVeO
KRaIhESJw09tQCopBv83KgnOkBp58OYRCYVjw1EU5COjzAGnrj7Udmy5GMwMAI+04gVkqrq5Oe2Y
I1ljTF+iAzho3A8SpQHdhxA/+2ZGmwYlQTwUVKDLlYRI8mWOetgPWupxbTV9GTEvzeMI0+O1nGZh
71Y5Fe+4tiqJW0xQTAsjviclezWU3kwhWi6kbz9gSocMLXHIEEWrOYcZ+xKXx+Bj/z1vWA+akgBf
e82IU4wtAgZLIYrJvcHAoUBQ5BeYiTod9U2DoEwDcgAwEwfVUDLMgq1cYMqENidPGg2XIePzBkVm
M129HC9eSxhrN6CIZwu0+UiQEc68RFs/B299Hfk2+fsGYiAUfdIkNK2ddAAslDEG+MuI8Ye82kkG
QhCHUlNgqj2XH/8PMma3XE7TpHcNq5tTaOZUoYjQkwZXgjwcHt3vj7BN87/67oNz0Y4k6fxqvRc8
x0uoaQssoCPkTkmo1cV9jYj33fhtul6lmIRk8Nnyc2nGtm4lbXxkof7Uuk0B2v7PJwqlv65K1lpL
tkOMWg/43fv+3EETazszDaF+jaNmckHrk/FxCekd6SgyGFVd1PLdJoZnoOLHVoIrj8ZSHSoJ3zPE
5wUoZjHNXJhmOSjRb7wO0XxTzwz2uOxn5/cH1ZCLz9jqGZnDEFVU3yn/pSO233xVu4cDPTWbHqBo
qYoZRPQ2lPufgcl+GXCcBwt0QGhsvzM7QAnMmCO+/6oQkkm4u/5XMV/61ZsBYmzsK22XMMxgMDci
GA5hObgz3+5kxpPgWnvFUfsXNNehGo9j7JwzKIJH4LdCtUeM62iog2wW8pJOtnMNq1JpbgPAISHV
CC1DA1nLHooieGIHqBKwEM6tbxXRv610SFiAMHXzFnABX5ORq/8T97lFeW10Je+8NJnYR2V11YfU
pnOft7HgQ2AokdXPkf0Rnj8UsxCDl3Z694tryO/re3FkLO33wDT3Sm8wtUudc8Je+sxQ7ibqiUcc
bpY1lby2zkUZRB8Qi5KsWPIby4tCK0EV+B62A0KjPakMxJVDph2j7LVNJE8ag7dV88DYERI9ZPUq
ticKW/TYq3bMSvAQgC3jxzDIH2NJpV7BINMEH4CCsG9Ta58QIFsFdFaAu+/V8WpEwcDJIcR0lert
htX8zGNE87TRhz5Z5MhgrigHscCiXi8Z7nIVZ87CzZsWBDE1VOzZ5PIQyGLdT9FLX2KGfJnR/R3H
7oZRH9BLAqcLqtLCxqJUmq0pj8j0mmjrp9F+ifKq2edNNiSxSu9HR3pO08g2CW+SL+1SbLJPyMdn
TqW4sRwLEUa/59sgi3ccHy2raZpqiSecscwM3SNEFr97dwTZS/V9233ZkNXtsLxGu9y2zetkAp/z
cByVt6F1XaJhERUgU4/ebfGCUz6KZ/0t/21kAMQkhHA57kPhDvdC2hwXdI7lxbgR85Gcu5+lFLxD
eqQee1yAuaCwptOOIbB7BSAcUPRXsWM8ZWnh5qXNpbYmFWpOpQ4VR4WRfuLBzSTx9B7yHwTJk/x9
mwCwNSv4YDOlVsqcraNwrh6rQKhaXZLBIooCpViLMTxYmHuM2DJK2uL+P5rpYQ6DApANMBVrnsYz
yxXdjCCQ2WG9oRWgwn4xg9Zrp98+7uKoQ2cxIYzqambG6+dXNb4BR5gDgSCg23ir0WzJZBLO2vM9
+++N6SICtfOm4d4lSr/dJ8a7CmYQMDO1mWQsLqPpBQHM4SzR6mvt0tIwR0VJr2bvZnkXMXQv+1DZ
iXgYVwyqphFsaHIro7VrsKC3udpWBIDvbhOKCpKd+ZFj2SjKRzJ2f7UczDzrjFpjvCFoQ/W1pWkX
nB/dLqD7dkmRKW3PLqzLVKCncMAlUodNO1fZyq1618I3O0yipYMjEwZRCLIqnGf1h/FKl0DRU9CY
JVqP+hETletAC5135oA0w1E6Lo5LR1+p2Im2iLFGdhCB5gG+smr6xigiKAyvQ14kprpRinxcLg53
cM6ZN6fHrBR52X8JM1gBI5B4j9knAisRJiWNLO4PWm5Xhim0T01WZTdXG0iuZ01fxbg0K1U52y1L
Go9oY/GtSWGRVkKvy/2z6Zgsp5ItqQHnB5CDUPhOyPH5sMcxoEZUM3Z/YpSOR3j0XXv+zW1XVoRs
OKrVa9LRfXz/TkMICGDfpuriPq+KfJM0+jz+MC45vF2Kn9m9Ref/vLYeYKUNOF84pZYhJ4r8pUOE
5GeQAZn8orGpUaRIUll87YrzgIv0N7cPp5d/R9m9LSHYgYDl8ENC76iWcT7lxSNlZKMI4+HU4PbT
qG1y9v1XiQDMCn09uGMN3Wgrthqf83U2NNFCSmnMYKHuUiSRXmUOANeI6dytWCrtzpL5Up1p87bY
uEvzMHanA++FX2LJSdQXSBU84q+9S/Iv9FC+DNH2zqY7lO+DKp22ClRJiaBa2O7FrXDZTVVj9sD5
e6PnBFVcCtOdE/ZdSttcDyGmOjRh9EhH6btxYfuljZRx0P3L0tlw1TQb21lwlLrwksahRhsbB0o5
f55ePw6sfCXb2TTF0WQ6hdgOnu3CuKPwuyL+6YriE6iG3UZDoB0mda95m0Xv0KeA/ZVjkJ7kkOlV
0rJfH8e4EzjBYm1wE9bBymSVX3RNo7UNLcrgj6xbzOuC05dGe5thAw9KlXpc57IIZ0w1sH2xGUhM
nV5AssZ5lANHONx7egZmefUp92HurSyjzaemRr5iE8IcUJqTz55GE2un7Ewt2OG5Pf6WOmxLrnq3
oGDpTNre3ydn/axL5Tg+hYhqB21DPor7GvkT3+gti3ZbVo89zxdbeGuzDCK0mhCW92t7sHw6fQSm
W/ZScfGVAeoAfslvRCfbo7iMrLgTGdGngQLF03Z92nInOEloh2IHksEc8ejjXuSnUUReI86Axcmw
48byp99gfwJe0/TyW01esHLbXivBTSqsOmhCKtoWJnhngHKMe5Eqd5twe7jHdsRJoB8doYR+g8Bx
YwdX3j821jfOokzIKF++jKDXt7A46QPAWn/gMZwG0AQ7A3ADzy7yTVEKhA41mC9yhdAhBwMw50dP
VOomY/XjtEa+vRVkqj5lFrJzuopxaNeum32iU1T32O6Npap6Pw3nSU0Iz0m0/806FxatvVZZeYm3
o789xexWd6fH5Dd82cku//GoOw4+bY3sCDYb7I+isFj+0wkinL8yzhyWw6N/5QJybbBQDK+9QTcS
QvEVBRKU+pX9CtqGp/eSjSur7ax2Yw08g0IcOnpvpr48sGp0DYW7lAsTCJW4Jc/vJWAzPqth1NrQ
Bc+6oFau1EzlFQ05kEZnAFb6IbQcbnDsAi/SoxOKRVUpuXEIgnlFdTPfxd97IH6JrHh9vLUcrkSf
0VAAL3/T+P8TbXHiskK/RZuFWX6q5eLLBNJaPH9mG88p3aMC5aPf2NLemfqVgsD/JE4moPs9LJw3
ggKxAzTr6sEn/Ll+WUkp5TEo7LqE8avfC67BeOnNiQEgXylAAXdE84PHa/24ZLGxchCrIOFonizb
KfwYry05YlPuBaQvzdEAiFlNlNuEEWuzq89PTEmN28YYKSiVK/J0mbe3K32TawK7ttGENZ8Hwktd
r4yqdISvx2TAuBYRGm2K8NbSBaKNyRv/4Gvs3KM0NNsP+7YlrYWAYh7Ru85BSfRHUqu+9x+9yLDt
o4u2ireE3uu4ghXBghpRADJqWesWyQOMBEFVtUp5Y9CnEMA2O0Js/g9/AzFFdNLCBzUqXUpHY+kT
hyMorY0zbpVulA2VOub/1dMyGzmy67NAqNWbYHr3+uwEzoP2pqCIIWvozDSRDoZ6ded7xnR/RGv3
1AhX5fdBzBfrQ1pR6buFbXAeCeU7v2FuZcTHzJCSOZ01tJNjPf7jJ1Ks8PjIGFP8mduTBPX34kRs
gPucUbXXFXzM203enz1ZdOnImyqiSw/FjNhAoXc9EnNU8xVwl2khpL6s/Hne7n24NTLgxwcNj8kK
8+5jcObpTowVtMqLoj0K/jAgwZcyMJuvVipFkJs2ZGnQAa2WXQQIVdhSSY49DHWsi/CgOSJrNHtM
IDmOp4Wk/P1dmA12qkn60gsN86z2gzBzyYLllveApiYmv0ROAWoCZ0Brarmh5caKM1e77rYjux3d
2RYxYwSKGWBSUgGo30pTLjODpJhx9QxGsIF2cZ1l4k5RUlSexGqqvhPSSBkIG32V41okpuLD4FMJ
976yQT5c6a9xo4hRaSO1K6gPCjIHVx3Y8mtalOhs6ueSIpyQ0lXhXWgLIkTu/7okTgLL1fcAw0NG
BDIzOwImJ9hD2Kze6kAQhtC1oBvezpZdpnhZYB3DgWFsYkGdoNieaNqybMaC+xPGP5YANnpUpH/I
VaSIngmdvkC/fO2RoQ1muRuZ3uf/KTbzlxSUvtSMb9cvW8sINEes16tA7zUOQRxk7fpTZBp4gspo
VTsxFB6L4ncL8NfKoVOFM09QJhqXdh1G1X77XxWpmvF7V3a6cDPG8KZwX1UQiUqdJAUhAApMz6mN
o2MeI5eb6/HIocWTgaNuyDb5eNS5doXi1y2QOls8EdTQq+esjfXHodXjrUH1HI1nkPjHD+mFTbuv
NvlagQuz9p4UXa3jwlpHTnBZzq7CJggKinehjzQV3N8Tcy+BtI+hIe3jPxDtpGpl7i9BqxO+4X2C
uHtmJqxxpAFk92Fi+CVYjgwpRQFPC6j43mXribwkHSJ4SUYrdEUgNhl4zubRp6abHjzHLGF7Uqfj
JcMWtEQVb9AI1QxaAIE9eR2IJ0Sj7J/bSjHOuPoDvK0DAhN4fdeKqjiPaMYFQv9uqCeUSUvUgZMl
6KMqouAgxD/rydBIfvC/IJiCZi6DDweTXYAbE+C+p4E7V8V8NO7ErEBR9yjMgqfY0fuebmzl1Tt7
MFB+3fTREUqiQepuOz2EYwmqaiuv5Yp8ZgbcreOxcXzh60PRty8khtL3s/ip/6wE/b+9zUArvvu1
YzzJ11f01i+OaHjdd97VkJjrJkTmt8HrBj2Q1M+jSgyV+Lxbp/i+UCyQTZbw7rL4II280Ur7rRnQ
HAs4VWFRDHgDU6dVkl0LlT1mdKLnmszQQH78DU1NIGyZN3idRxhmpXur8HQPUbhrqtxXwAO4jmBR
wJ/Aut53vOLhRLm6idep3RcJjMghUQcEFEa723g6wzEc1sAcHCb6/zO7fxMEb9sZSgd9OIG3DHwy
lTJ0uq3yhawtT9msZrtMPrX5xWgJHoqSTJDxNBxSohghavvB5YK4GeEj0y1uWC6UP+S9smnNNWaa
le3VWlGGEiZa83xiBS1qK0YUUlmNemdxTEyT1EFOHvVHYgNuLE0Cc+Yb9j707Doe5lQf3m2to//j
ZTYL+PJlLEHKHujP8Sk4fI3wnwKJPUkYmL4iAx7pgK5PAcGrm7leMmBB28YbFEE16cmhKuc1ZAOi
xaF/1St3cfWPIB+Szr9yyEw+R5m4L2sUwLGI+fbF3Sv1NJjZG//4aipZ+Ygx5pFwF8eJuapjYpjL
J+ooE9wy5lnkcahuVMyOE+t+nKNKlYv40MAHLf0R85vI48pDDLRCCaA4ZHy05TQ1qRuQf5WxRY+E
uXhbMpBOiGtJBmDAm/e1bFqwV3ZrcSMj4bdgdND0Y1RtNnoO+Y6u0SRbIbz4PzuvZDlQhLKGWNVZ
30AeO88bBzrYO/0YgAl9sw9unoJ+7Zgn9ZNVrAhQ7N+2FzjTFCuI077C0ZMMGvwpjX7xjoTv2IwU
8Df1hbzRonKmI4pzkq/eGkOfiiL4KWSMtoLCWiahu3QJLxca/TcRM5jog7mUAmUv4gEEpBUh5eak
fvaBOG3uBctEP/7cYEkqzlncux/uRoeTDwRz4S63CoAcrFHru3Z3DK3/lxrofaGU66rzK78nvBXb
0fy43gW3R3xvAcKxo819PXzf5gbPA3J0yBrbViinci4gGigBCkDlswdkIvyMe0QZ8iKRJONh0a+/
GbOdBBbi3MCcSVIBP4PIffqSI0MRY4/iH3mt09ujkgVw32Z94RPEhv0RHvEpo7TW4kSlIZG6zXAH
VboxGxMXUbsCr7A0BnhWLtdnUVJUwKiUqdsQddxXP2dXFWCgcW25d1bDfyhK61IELmWlMP+NGLtY
SdPJYUDIC1dYkD3k9BF5PIIP1gEn5nyIPLoCEhnvAB53t9mLgb8xs0SwELSovl8iOxPohWgbN8E6
uHnEmGkjb2cpySOk39+2JS1hZbJSBNKDfjc+hYdj8xIAy8Kxt//7aLHicbQObEZ0V26g1LqHTiId
PRtq4yJNw9nR0VZ4vfVaHZvOFmYBA2WDJw3zLA5mVFiQZ2lOprL/NDKrSKGZIwAB8iB2Z3B4RrhE
L5MHGrb6D0115SUszHwyhlVg923UKwJVEFn9M/6kYW3jBsjNMEBnWb23oB7E/1bL09+hNRqoTbvl
a5swctB/3QvVVD090ytHtnlSHZ7HvU3CINB5sVTrbrUcF3x9SEWTHseVVwzyndOP0eC4Kco5wisp
nY+t6wLcyms2ax4d/yoP7YcOshrD0V+8Qb41pOjSdY00OiFt1N+pUSkwv/BEU4EbEZhrKAvatWIY
iQdwVJTizCmHW+uqklKfFSHL9uAAfAAs+NRWSm2Dwd8BinFTI8BXm35l36snMUwlx0AZv25aQk0J
qpjYzsTn9dQFSsI26Os+8Wku8d6GrcXBRDgAJWT1/Js/uxxmyQgrjhndi0MfSnGKz+N8CNzmdHMZ
AA+PYuYH2la0kPjtd/JQztEW366IiDFeCmwYE7WRoxPyj3enLkmUg5e3m285/JJbeikeuWqXrQ1h
xyw5ls5hNCUeh86qXZK2fwPjoV/PiPe4ChPxczTY4QKDCsX2e76AAZRePqCnK6P84XyqrlfYgTQO
CQYVzybp0bBWMGCo0obaQd0ushlinlmVfYAVcarRg28USwE9kmlVXj6ZRCC6XmaBIM+LLKNZIXg1
KMzgbeMoId6eZHn9iyXthku+KCfuK++9gFlKWeBQBs1fsf7m1++4jh8xxhKJFj7x8wKDHpcJ4pNg
tF3qvryd/DCyy3pojdju/tkP6bIq/YgrlLS6MGwgAko6mmDXMf3E/Bm/nm/1lTQu2qbQfxF2Jka1
dRNDPEblBKd8nmGTXCnc6PGSSDneImkUzWOyATwre66EeCK6RnQM9ImdWKTBdGjdIqMez+dTGYcZ
N17Ju4LcqdqT5PhwKLhwYlKIagzQIS3UcFDPD0dmTxDlQQM8+Zy7B5ZTr9i1odO2pfPEsYYpRrci
Q9bIq9XauhQF17vdVRSPRHPcjYqltHN03TmHxjgnJmyh3a+Eho1v6+8Eh60+rpJBQQP1b9ogFtUJ
IDNA0P/bDG0N2ITJNRFtUnjmcsbifsj9u+HROB4U9e7vmIWVJmxIl40orFnsIxegHdBJqHQHB7pA
P+A5UspLbC+UAZXTzFPOeGbiWJu9ASjECALPYsQAFDK6FLdgzF+nir1NZLhHdioFibEkuMPgAMBJ
jvwFCSGmrzVfQaWtjC09ATUn/+r++FFWbBu9/Awe+WWRU87IuKuaTrsllBgT6P3rMFaFGbyjutWF
ffxbQ7+9dzGp8LjX6Edll0jA8p7oHySCeES0uI49pVVkFy2v+yq8reIRl/rxaGg5+IJKjn/3uF/3
DhI1Ln4hTcqCvOq6JG+wgaOlYoe/ZavvSaGSw6jrRbGq2zFAbFARfH+cfBXp5coAZq3mdX/+/JP6
1PEvLHTXLx9qXOTFQrtQ9QZqNC7pggfKKMW0aRgcWK4sxTU5Tur8Je/Gevte79j4MUAbgqG2ES9a
0JXqqr85/dh0aSuFJlXaVjKHsEQzPF3eeEitlXDXtdRl0Tzpt1gW2fRshbaUYCKQQHHY0byz+eow
gtx5yMB2dUgpy/5e0Rdghfhu8jnc4CwAoIRw7K2Avk29FB4LUNd1FJBadBsmaYbx3WvQW386fMro
swVeqCiRCm8S0wHAjxQXonZFE8nxchHbjwmUcKB1b0yyzwipk1U5TlVwKgbc3Vi9wo6tIglF2ixx
RwA4zUMlm6jxwDTbfC+P4BkFHNnDS2RRAAk3IbMfCPeaqe0aD978c69CmgGdO4BQnCb8rKxXAdGX
lwvg6A9j83Hw6an34+dzwyzlYtpE53cQ+BzYzX6SrryJQIQEimGgtHAx9mzHIXgxK5kF9T2ox9S9
QCYYW6AG7/QR7/PpW11Vq6VD4k9lmyqvYeL94M3mmwkpAEz33zaJAL+WkdjdOWFPehG34Yss8vZ0
9HPGyjNjUO6bTDYPFlufm7KNTIfXamY8gdhEX/2egQ4jLb05PHGVzgRW9wgDD8QudUJI/MWX0mXi
1H5sJSkDdKC6jSsrVxRj9KTcmOSryYd9L2dmlvNgYoryj1c50I/JFJPHBPHZAr2u6HWGXj6y9sLq
cvnXNCKXTjBz7LCLN0/LYKu5kDBAS+kAnd5nJY/0jICovvJL20iXyqOyCz+j4O3JWWTkWOqte7n7
ixN17VPSFq41B9V0gcE541IsEKd0dr6x3HYTV5l+Bqo89fQK02D0ufUAIj6BQtLfeuZtoQcsUIez
OS/jVlu7/Ooy2W2Y43+76i37nzHJPT1FEINCQZE36CUUf6+Pi338nrh3b0Vk9J/Ajq7YOmm2P4uX
p2VpB9L+4SDOneydKaIqbVyCUBuitb1mOjf75HW6xeVxIxnZfa4vWpSjDgeMxTGtJfDrTYJULhqu
ibMJ2gfh9xwCzRoqbxoswYX60dSGEDNlwH5qJEWdXVzxTG2FmW2zhw0hNLwTDWT5NDNarOsx0/5D
2vGpjRqv8H2vGKRl+TxZFzhflnwxNzyq77veUV0AiPkRQUd9gJXLruKZQzVjCjSEp/M8oRr8rIPk
rUhZVNCshi0waNouAexLIhmkJu0XL3BcbBLCsjh+NcMdcFQfJZ4EG9rowovyKjompGxVSPdAEera
mvMGzYpUsFyCvU1Sm3P1KLSxmJdEC8hFN1I2qgHO5nypSZr8RyesNyj7+og/5PeuCE9LCjVK0Zi9
PZ3s//HjXqA3c37uH97BxvT96In/vaBjnNLMjfvyBk5uTwv1IufLncRGRlYDW214T0UaKJPaZJ9g
9ZWsIeEXk7l0bQOdMSwnHURTY9ZpNgHAXoa4F/J+Dd6BDJ64eLa1aToGLPsDg95Exkn8nM2ghv6k
T5hSA0jDQ6rszyZ6+7FtdB4n//4fAyhYEK9zC8AKNQSHWKW9tA5gBVl1Utsy8KmlefBy6Hmv0tSf
R5lVLYRpqdeR7wNmaj9bH186WLaUBPih2e+hDzDuGof0TRvD6TCWUCVOxvBx/4YVzoTJJ0QklKtD
mCDOo8gfgntmlaAMamjPZmeLcdkiWG6+mOBsRoQpLibbYGDdinkwDv6+yMrFQUegS/DHjb0135KY
4MZMYf1xKVM583c9Ac9hFK3BuBt7Xz8+kPXexa4gcJzZwgk8Rs2z4uFfIZOwQZYVPQRvkTQDOO0t
3xsjofwrnLF/XKnpbcfYL6q8tJnwJHiIShHReiWN7MoJupDflcIpxo39p7cZ+h7ayvmPW+bMw+kh
2kvvQRf7ipSFmunP5ZSdIufu6I1AR1dav+BU6KqT/lQDLCpJMBydY5Tik0Kg5PkqNxtW+jgbzkLy
kwdT2/Gfhw/wmMXIdBfweQVBzW4pQX7Bcz1EqGW2jfJ8c5sGBAypxFzrMkP2gomcO6pZBS5z1S7o
0X5gUruBJ5KH0Q0lrnXE3hoBaZBqR6UaB9Pk4oHi51+mwk3FZls3slal7VhICp8rVYX3MNNXCZFt
A0nBTh6cvt59czx741PECVnSF4+kMv8Cwe7d/MT9eQcvj/e97VgLZWw33tVqzpoHxgn/ZAjMtmMH
A5/TF3M9IWlF1c016R2OLB4UqyAt0xsYfScnI1j3ZSSjOytpLr4bIlNT5wLVXe3Ri0HYqpoWf/Zv
PHwkbwCqums6wcVqJINiW1Ww9LhOCQjEUGYqiRJeTZvb9lvDCwoIkmT3fYff/0drCYGQdP3DQFN/
GZEgb+K6HDaj0dko+P31bgnSz1XwFK/M6FRwI26SZMgoY4e/bi4ODNz9fhXaLlJRIBVRMhn+eh7Q
SVK0ydFr9V2rPNvGc91pfIV//dAq04WzQi28J9Aoyv9J3McZIDwYCOkaAfM5OsoBPiwTTHxyrTJB
N1yLHCclwLMGYkuqpFZAPhLYbB/jwPoPuAw3PfFr9k1Fx3aeoGMUQ6BA+QmnqN4NCNaukiFtFttF
oAMc8eWLSFHUd6OEFW4/U7LmTQSXGZSKb3qcwwUQAUgpQrBcCMtlBfEd3q6lUEDOFpnR/1W3vE4S
28N+S1yVWc4DDLiuPFvdI7eyaKP/oY+AQ+YpMmTMB1d4PsOy3zBp9dc7+vf+pqFcPLkuA5//HqWC
XZfnyURrSpj1BQMYmx9JmvywHNcKlX969+Ri1zy3JyzJuKsVImSJLTIifbUJA4BCl3gRbdhLB6us
q+QYrqV4YaZ8bB8jfstwsEtwWHGovTcALvp2ohHtHFO9QCBHX0aP3zTFlYR9M2skKO0S6Isuxm00
91pWIFzH2H7pbcY86+9Zk4hBnBw7qo1LkHIoMljONlDcd1ctet68eeSuLBqn6eNMA8pMniTgtlHv
EAkMgZmmywAnqhvu5ecJOAn62oGq6bHmT4qGRncW+6Kqp0YZKJ2pP1J3nnYB7PkjkTiBk6eJtahv
M+AyEz2llDCbw0e95w4TRxCq7G48rHE4Ty759Bm5CgDugH+y9JHoncFtZlekPN6RrlDVle+IUHJc
lm/T10MCTJgEp9CZ4ewaqKIKEF/4xpgBEyXQqAhUU3H6sbmK5cErp4QeOG9/QAue5fPehWF43ZIR
WccWgeGhnHQyNhd4jOv30+QbA5lMIx5imJ5C+/2htLY600riaA3SxuvnhQAhUgufIPGRsY17vph9
BgHySTe6vzKhRsgFH0F19AfJ6cpLuwrVezZuRPMv0ku21hNR5Z3fSGYp4tHW3n7gZNn5VJM8AqI2
C/Y6RFcjVC/Np+jSR7zckwyKJuzpDXG5qcggNeuG8AhGYANDiNINgbLMJWusjLxbj4aSlkKJpR0q
uvIl+5s1rEphywLYUXuCAuTZnmfd51AYoEk15yFq8xoQORToyFwGZOGCy+Cc24A6duwm27mUTs5s
3RMRyLj3fPAEH4Iq0GaNbfYicJc2XHtsyqVyZ7coIIipvHA4xsJeUaRNq1W6z/7/wO9ncMshnH53
jzRm3jlti9iWzE+NqGKYR6HZ1pvPZYw+A46S77iWrxFeKQzG0P9hATFwVs2tfmE2UQXHqJKkcVfU
9TbAcYDuCFaRE54FSuQJq0h6M+BFrk1lGQRcpce6x95puI4XwQFUlro6Ra4wlLfMvQEBlj+Wv5s1
WCfiXXM9ds1hyk8JP4N0Xu5kKeKpO32t7dIWTWnWBjoP9eZK+MmI6Y6EoZMCSKpyiGvY8G70l3fi
/mpYfTn2oHBOF7vO64p3akDDuN010WNBXY4cP4IRuuL67RmqPFUVCtTPnleZq62QKguLME5JwNFa
0hqnCBNQze5CM9T/ppVsJ1CLH42zn9zeNh5d03AFwcteK4Lssdt/7ykXpSLHKTK9aVCMsqwIAS86
wx+6HZ9GgDLKzqMvZgapfZWesO7R8T0jyOU63HqZnsJtbD0JRzZjrLzOfpUUGZMZQBbz+BOrMdEm
We3wIFcMtuF++I65LTQoCvwEZWTxDhQT0DXO1//wUXX/wZqdSQ7ClSoZJpGYbk4X774hU6H7u2My
X/lFyKaLcaC5jZALb/WJzTv+4+ph0a+JUcXI3zUbCjDAfQb0NZJj8KNo0cTeApvGSTr0WlHhWKcU
31aOPMBwobtl6F+qyjxCxelhkSPKH+9UchFjdko+Bt2lysvu5P4G3/E0fFwBCIsvGbLj4p8iz6vn
vXR6wbliXlXP9gcVDLpodEAceSL/ri5R97Om6hgngZRR0V8XjzLsvO5EBuLccbJLixd3fRdQEH67
xADZU3DsV0q6f0ApBPbLtH64pPTf+7bdJ44Qfi3lZqxMHHpODhS3w4ugbDO5FlTF/t8oXjtTH6Kx
lWIB9KTnXsymZJYqoHLiDz9Jstuj/tb1H7DReesmHiOj98xcCyR02f9Pzra7oUE9KCFoENmFNQEZ
L/ea7psH4/udmTXc87EYgVk9r5xhk4tfdFqgq6Z4HMB/F5UZ96cTKaRLTsLDdZKXZL4oASFkzVvV
wViF01C9sAv2A/Lty/QeqcMnfaqmF57ba12DmiYoXxVm+kzWGIiyjgEvskKsVBHa0Q8slC7iy0ui
25K+v6XgeEZLjM2X7vYfWKcicyom+6Gfpum0gxErhwo/RyGjM1TjzDuTH/O0sF5UqSZ+hH/bViqz
r1b3uFLsK0fy/bcbMNXE21Dpgzag4SlSkDXY0H+Lo1Uci2jx6Mm6JSXyRQ0/6fl7RU27qourVaFu
UyOHDCbCGNgG/vEB5kkEcHSYFx08sFoGp3kGjCc0vpTGOsj17OXEpALujLj0nxJhN9XwPaZ7+6hj
dtGW+xdGpMtpDRZPjt9LqZfoo3kNnq5Csy+KrM6KdCUkQRIzPg8Z8ymX8Ei4gE9as+szJpAUbVyk
UjpPapnHTek3UsVMYex7xRnKNZfZFVjxU3BVVbJVJhHsR+4hjLJFmqGJJAWW/OsPjuqVUknnk9uF
2UcMr7xcizcbCz6XYQ8H+ddz2XZtWV0DFS81wf0yLRrnx132CACUG6dK8Yee+iaSI6wd7HeQcqrT
K0LWMa4YxTwBafscOIkJGqk75QiFPLHIXIfSODGAn8/b9V98YfljPd0vjnEhxYioZDkMQF1nl+zN
HDRBUptvMoMbw+wRlAxnBe8CdnGc6RV/xlRrGb/h2T/hZeFw7GQ0pL8mggtMT7m4QFWNv1lRj26f
dIinX722rpQSzBQfBHvVLXRuDYhZTCYvmiHIETlIf8lpDcW4CxB2ndHkGpb6srdHKtrCN2eYjbBA
SREKa2WUw7Yq0fFbkmXXo5yNLz7KpYr+XhuoGXLZguE6Il3WD4KlZMI/5g4Q1K0LKgxLL/0KnZmL
qk7X2BJhw0G5lii/HFvPtKduIqthwKegPeJmfq2/em6gIKODHIZvgi27ka673xoQKCUAjAFkcX7Q
Ted2A63ASYPRqa3kxRC9img4lXchzqmgV+0z0vGoDFeY5k+bI6Kpjt5ZGzt2k9bObuwOfxgmV3sN
KbVWCresrek1rryq5+XBKwriqouBERsjZ2jdZoWBzG07jif2jOYg0m0L81farahVMGRMOgfYc6rC
r3kOLxAMCb9Xnqu97jVdVUOz9+OVOqIB0siJhpyh1ZFS64SaFKZ8FAoKDbTyj2Ab3yBmNCUM63WR
7Z8z0qWG0VyEw0XEka9IC+o8L/EHotcM+tCEY6cQh7w/vd28hdT6mKSUfTcKgwZwu4E60lGVLzKJ
oee2081geS9RWfVRixgFJnNpaFQewnZ2yhnDDC+GZK2pbRDJdtwNHN/wAy8Dk7/8JleeSNxC5hbR
mc4ewHQXg+Fncbk6XNjDeAl/MQU6FsHrCWF/E1dP+ajg9t7bdRJS/EsavJKMSX2xdx7r5q6S3dB4
PBHbgEZLi5xOhNH+St56GUCOlmZk6fkwfaCiTkwunkOW2fTai29TA6dXIzbZ4ahQ8t27lTc+Gvp1
W1YCq0r1Dj+2XF1YMRmuJDexyWpQIbASZK3Ot7EjsrHAxF4IFKr4bovzR9KmI2X3qrpYMtUvZrby
lCf/OjbbeFYS7mc+bdRye/LyWNcAkj62YBomIQ8X31ipyYVu4OUpTrNJIQ586k5hmiWX81p9CkWk
ZjSCITZLk7d+dKR6iNBJridOKW/mKnETAd4xIvU/AdIxC+ZIwu4newG/EbfdG3v/g11PYV0x5XzV
pJpaoR68aJFPjJpXgXVyFCv2jU91iSnZB7q4yInBi13o2ckLEOPWuF3TFjMkJSrrFA2UZw3Ifduo
mffkNmXt9LwU6KJU/XPOovk5yr04sYxf453CAi09tgHCjkZTLOu57kJzi14LiQoKIeWRf+lsemRz
l4xSutZSS7bgB20MF9Kkpb7hXi2TC+Luoz1CDnx1ozznWZ942pvkWA/HgwAQ3k4auYSw1vJXKuBx
PjPWUYx89O2LozyL7yD0unX93YKLQjYSAzOV0mf+T3gHGWB1/+g1Ai4EseW0U7Uf3Kb95gOXnI7R
IdpgI0hW3yEahJ+RF3rfefRjbJRk2Iby2E6DVkASR4W+Ajn/FhIyqlcp1vB5YsxO9jw+kr6XR2Ke
zFZZ6qvwmEMrs4WAkPprZlHxs6SEWt3DzD0nQ+IDcsJ/NSW3Dg8OghQoyBDbotApMqWOHKX0f6xZ
VXekcqx5/JO2okFNKt3vZ0vzEYQwhodb+gkwWD0raJsvaqjjQksat1Sjf1MrK3aT3JWo+haFX2+k
4OscewvoOF6ZXi8oTjHpZvK4ItnmaWmJOXJDchnXwtuwJPkKUc3OmV4JX7fRnbyTG7kxdNYOYwsp
9rvFXYo7/+z7ugC9xW8kZy4nCDaAJysCiNh0POuTL3F5BNv35GYI4h3fVmiIg1U0NHYOQm7N0nHY
gRjwo5VtX1UNfvhBQa7UoTJ25z1RFwW8fvRwR8xxUqKIvd5pxhk7KP2Ua2p+gQM5eXL1FtO1ubVy
I2nQvuZpkmnDHzeJoXICdGozXnJA1M8oTSf4YqicXgibFNuOE3Mm7GQLSxQKINJ3GNYNqh5DK1DF
NAMFbWDp6qpygs4x3uCUL3cYnNejIfFAyT3uaWcVFgn5va7Yq3VYOItgVCiGr84DEPC6cOyeabMD
W+WrPL9US4lyobzRoLzajdDX07UUffKffIXRpUvnsxnyrIzJOYF+QdOOwa9m5cpoxMQuA0WqU2ia
LIa+6yOK245LHwIvemkZy64U3Ft6f3JdY9BmfYwBjx4UjdvrCqJXQ5+/PitFtkAm9hDVCd+mP+QW
Vh3c5kEFFqjOmGktadocfEXgicqwmTXEwlEo2v6od148V/VI79RAJinIoO7idslwJSJCdI39a4v3
f/oy2IenlcRgLVVouQStiTRoFv5K5xSRDQWRWmvpG1D9koPZe8c7oDQqm+l+DAaSUgnCSdHe8H3u
igJMxpWS0bN5luuoS2SErNaEj0AUqQtEnPCHKPCCIsRhv7Rx7qFYuemv/A9DREdUcjMTTsDUNxHK
c/savNYSOq++9vVE9OgPo+MbKOPpgWegyZKKhR2Bt3ifOfHR/Q0sbdKWwUWmrrK3awY/DhKbqYa5
hOym9djro4mwm5uXEEwU+kuOgJ7CsSc80gK0nyI3W+FzeY6s67HFb2MmLukUL59xHX9gohhl6dJG
PEjzZgDfKqhjIGa9kEDbaACVPxxbhuc5ZQkvgVtFtSeYs1S6dKIosG/uXhdRB0M9UoW9twm0CL8O
MKe3DXd7cA1agGQoAWa/gYbLjlmCblY/Y50O8CrqFgxgtObj7yTbRh8Gg7T9PaDp4QmvHPj4jhGr
d7V66fb4bPMIdfNSQUGw3w1eBcV90MCO8xbUhWyZrNaOmiSrUksM6UVXZT9XfsZ3WbZ/qWqY//sy
YiNYwPijdKRddj3ZpU7RQD/Jcp0oJB0NcXGSAbd/I7/YVPF/q0qDdjqgCe4WRZc7NZhkk3jnY8lA
nJoC1XdlOSM8cSumo32WRbRRC1JgYOXwVtYbfSZmN2RjUFdO0uZBhXiNoEecHZ8etowcOuk40yb+
RUUOM+YRODpCL2G7NN22eQQVcMGImdzTH91sG9jrK8eF1roY3AL+zTqJMno2J85jIcCZkyUZ4GeD
J/MTwW9EFmAvEL9s7Vg6UHsbclZX6Ulq4go1GHThQnQLZcx1axDYlGyWV1ovkjKylxNn5rXhKhlE
yg81jo8lDjGdFln3QDbiLXnyGg3Nb8cSRt1OfE0lV9LLYYNvCeIV27FqxiKJaHCSDhYcqrp/DX15
Ny3UtVbd6AX/qI3e2PrIvZdL//HESmop8cQuMHgd0M9O03eHjWGqJvea2YsCi2qopdcilB1JihTh
aPjjHVUB/Ssz8rLl2aiZEdnwmqo1XuJ37FUGgjf7B7qTv7x4frnUeuuGzPnrBd50yiWb1+6JGuWL
o92z/1PWx1vWYyUz+owBvyGJjdT01U4R8eTe+ZLtoTEB210SXQ5LSadLtRuEXT657B+MSWl/wJtm
ZG8BOKRyCEFwwgn2wiYqcMSLdKSxYJFP+43ZfZF0XA/YdwpygBmVRbuIzVbbDfahZMKQnWJQz897
0f7QZZ3FB1PS8OSdRsb0zbWfVTE4cx3/+QsfEWKFeuxBkik3a/0A6aLnq0mvXOGzkBJFTcFIP5hF
nxhI5TzeMyl3lIlB0Dr+VOWmbpwv29tmvg77T7KPEzuvl93fN0D1FS6EJD3u89zMaZB0Rpy4ws7E
aQjKacy5zj6fqeVPyB4+r0xkmz8optS+KHo6Y2VkTynBvyEwdt+eDfwHUMmcQk0YOONPg5LOOv5G
dr97k7I0ja7p2+h1E3LXtcfHyOJ4o6g62Uf4k+GDPIIDjF0H8cN3sQXYSbYK7+eU6vLvfNpocgTS
uW3LRMev0hDsB8fx2NnQ3UQVzEL3Yu+tgo9m0zY9evsktQDLjxt+EEcU9OV2W9BPSbA4LJSdjtHB
h0lbDpzJlnFx6jDJz0WuA/q8HQq7mnaLadvnShKba0rce/UkdVEjF2Xx7k6XqeJqHPDIhho3fNM/
fkDeZ+GeqCX0YuBIqZPKyKnoApJirY/cjR1sFWbk33xZOYrgMj/oC5cCU2tgXoBakDAVXqgMKVMC
PQ3a6dyet25rm8NZIAlBQDyJ+lp0gFOOxG89sp/1sYjTkKcHUqwI+6wn0DCTVMS0KRaSNXH1SHpX
S3neAH3p38qKn8Peec0hAl+SICWa22rKLYjWxsjD4z/zzMm7lK1pv3IXD9+cBySIXNc1trv/OwIX
iFOjEGvKVn/OHxELAtbSs2lK0uPt/jTsFa8ajkVaRMXsHxN2ACWEDwi4h3JToPaeNP7am+e1Xtx8
StFa3RDYH23XObVTIMKn+OIoAODKMhkzirIkwWVQqaTbFmbyJ1eAmfsyNWec1y1C3dBKluXQl8L4
L/3hG3F0bimqYcDXYRgxvIeQvHzwLYyKLjA4tVi8kKvLu8TRZ+FwBI8veeJQCuo3q9rYnGqkkPAt
CaEGuseq3nV+ityCGgIQwSuWf+J8VmvivBgmofVV5koRqEn3ycbG9sGaWky59TxNyaOo68Zw3cw9
YakVPF+f3kEcdqrxspVijPImRBE7SA3sk99WrSLrFbjMWGvFFqSCcXalB0DZyA4dixV3mzdd5XNf
97hJ0R71qR7Aqdq74uwTtbkeWg/EkFKubbUs5Hd546V+QCZNYCE3a7YA8zhrYq09V/yTfKk7a5/1
Tz1EQFJElvb/0ZL/PpcizwGc2uRCMRWn4z+CJx/I+nz8c7YqBQRKUwNQ6FFj7zPuz17e+VTKeKBJ
sBN+/eCL2F+/p69jYrqZjaq47zPt31WLa8WxhhBrIJ40ib84UeOxyz9eGc+RrrmEhxSafHQvRNkE
hFyRMG5mPucHrxZbdpUrZuLbLtYivCi9/T5M0I2mhGkKAGm7uZFOtyj4ZELhirdbimG/DEB7ObMi
iZxL+wSswu8VMCvKI/Fl/czIHZPSt/w+c3YUuW/I9BGNeO8KyD1dMtLWCooQ0IoxkalhpTyYwB7z
iz64zBUWmem/VJh36ui3MKV3Nm3xn+DLeQ0ZOUFBEI/nt9Epd5n+ot+GhIFDj2alMrpIlXla+jlS
l+Pd7fC+BRFPrhh6T+wWCMPZo9JeB4ic5uVyvNJ2sSYzl71fxPjUvpWH581oWAyofGSUgIxnHJJZ
xM3JgugStS6w0M2/HBpiqzxj+7OcRG6um6KQtPB+RAJK8GdJcFYKLuK13rkLzFlTq6w6eY4Cq4aX
E8WVzVIeVGEGhATrq37/Dg+hvLEwFPfqUcZC5ge83biX1lApwMd81DUXRUQoPTvJms0P31gdGxP/
Gr50cdBmOekchnbe3bEKArfmTbiPGw5hYgp4sX1AcOucf8x7/cXOWTKE0DIcHolUKUybDCEHGYvN
BojC5Son+1rhgZch9bHugFUmtWUQ5HT7h2BFFsIOTFI18qD89okghueS/lZd0uqAerAMujMly21M
Ut1vZTubfLa4nQmcyeyts6He4HCbaNBHJeZm3LOJS8Ip52Wbwugeu/jnzlg0FQh95kgmWjRyTk1g
MDE3bCAJbHRRH36q29AIcNKui+40/ih0tLvi4PryatLGipk6DNyCdTW7gLYD8fot0LtLeyo7nzF1
ceiL+6DzSVTlo4dOB/PGxWriBlfh7ii8qTD/Pdaw3ThHed5iGDEe1LodL/QRrTanNBSg/mNSeWLt
jlC8sWz8MWWM61XMCxfOn4JECpoMAiAlu+Sg8E+skqykouQDebnRcQcCUxnThtZ4qJULnnQb9Osi
pziNYCZIca9sPbT71eaKp/v+BpfH8M+Kt86t+W/7UlijOzkf+glM56HrQA5gnuSKobjhLpYAqpV8
1f+im4sFGF2anNW/pIZVErrMd+j2OygiKisKWtGdqdoE1aYbjMsvnXjroDgIc/KYV5DBjjWDXNCr
eSwXUfZRKtpMAED54Xr1tw/FhdMc5+INmXyEC0wts0iFoGOOUmL9ElNoHIdsftzB34f9CJTGA0RM
ojq+zPtt7f2qPb4o12vCKWVj2r1K2QopZho6yix6SHMMTHru641xoNX33WtDvPUWJQef0UeOsitx
VpRY14seaxpDpRyM+tNxaUHtrNFhI0tT+3/JXtvkCqhvGxyOgBBu8wfXffQfYMWUD6MvLwRNs3fH
cofFZkKerLZlQ1vPDzsPDaX7VtrSTYwQ5muzWI4ci3NR+jWHv0TeGgQFd1c88Y3/IFcbXI6ZcaE2
twITs2oZAN4kgZnAF40Y6FYFAVAh/IJ6fDVeAHxMXU9NsKA47TzZBguO31W3ui7WH9kIdDA58b8d
IRlA3dRlo7Zd2NCHCE9yA8xpm28FU4dyd/ZPbXr5YUQl6swiS3/mlLObE6GpM8hu4eGZbL9t7Rbk
/yiYVhy90bbvvwTU4FoPEwKop3++usNHb4aHs7QNI6usv/WXkEJ3IFODAhw7m87OVA7IYsxVZyNn
xrj5dQPvKw6EGrjr0XiNi9HesDNZ4Y76pw3ZTU2kSlxXHwZ7N1KqWYih5KJYkHORmiBi5Doludr/
GLKTuRP+YmJckGUU6u0X38tqLh4O0REGTZMFOKOBhCqi1cwS64Ty7KxQqwylUXR/IXON2oAQZ3g5
Qd9nBlDr54ziU74O8d0wMq3JI8mhTOAadVaEV485Prf9nsnVMGVYUjwwc/7/yY96DNJW70suZEM9
/umSWFj75h280qBGR6f5fbW0dAlc1SYxE6RqNCBrpOp74OB4HSaNyQ62r9KiXRQJp49pAAKHDrL6
qFtKyw3T+TJ/Q5wBh1+wOxIxBiXRVy5sejlq2mW43Q+cTXQnB/Pah+yMW6x5sL4iU+hf+NXSWLz/
D31YKIEs8Cxdyql/oWKTir9g29WnFIg29LCZbuQsA6bnZ5/sNgwi6OT3vUbJxcxt+fmZLN3jBlRz
ykIir8LE7aC9EmqmyBcYzThFKwOQO8d3bI7djAqaqWH4wdpkRtXSANPzqeQTIiko9MilcHQPgNnx
4Tp3erfJfMLez615u/GtyyDC5xkUNokVKNUhjHrUfXmTl3xkxDDQQufYtqgL/oI19YfcfEn8djeD
qrcS5OllHFdFdb08qKrU4fZf8ddvHsgD8VUr5jkAI3YnN/WC67cEKJmrEKGBXvL3fdoav1PG224D
7ORizVdZ1tMFpPMZJjwUmvQ3KolPS9ZgbBo+w9AlgOya1ECJHskeiVkEfKavQ0PuYFEBCXQYkuio
PxIZU75QrOVFroM1JZoMbDFeSNWjk/1L4jlT2msYcEqM4wjfWuiTf7FPOG2yAZkAV7T9bxj13v76
oz6WKnjMvTX6YDA0ppyiMuLuit2Elw4WHeDYflJsPrn32i4qd3XIpYDh2HPjCw+eLulEjes1wZeY
0gqJCkAnRKwZSEwOAuu5CP/NmAfFaqxBZUW+7F3qFhQbGdFYL83HsoEb/aqccS33bQXCbhed6GLw
UTZHpXeQqOHC8J1JJazXZ6Q+q1br3poLkpfnmIRPJ4SWradaTtNftLLG8cTarso0IJr43wfMA/SQ
h3DiZU7RVvD4OiW6/bpbPwWEyM+FVGGUVY05UBifISEMHMTrSW3S/s2pjVfRssNgtJ4HvJDvXPis
bBAYCOVXX9W4aAFnsUa+JZa3KVQ8lUF63+Y/XgBYGqUPsoJb526PYvRAhTYHQDi65VHSjJe5EILd
wcxS86Vdz7d+Z9hvx0Dz+ROz6U0mo9s3Fn2SJ/Zn4OaLWVl6UirMs+SY90DZUXV6+rJyibUIYHCG
PhJgIRUPoXNd1JuZpUt4BdD0BOvwmVRRClhRImRb43unuE2GkngXvI6dcYx4fHbvvXp5O0s5/iDS
HktsvotiBp+Cs0PKDcehCbvvvQs0k9Gun+uzo6ONhuTtGat01HWKJmlv3t+NgZ6OC6nTv0WAtl8K
HRjGIIj/Oo6VOkTO0RuHFaXthzKgou8J5GfmiUG5z++4NZL2QyrkEV331AnLwIZm+l9Euo2WX8q1
1peqZMs0/5r6keoIk/aS5BsWQUoycVA9hkb2sVePnsRMqNp3B0Q3IQQMaY2PqoeRyKGUXD4xoHhs
Tz/O4fX7vEMpiwY+mumDL6owzd0pMEBJ3YgY718IclXWJTp/zW+3mvir6K+einh6Cpvszz9dvrxo
rkvlfHgFsvO8RzgrVglCktO8aLzZCSlTcxPVM5WGKScOIOqs7VwYwoCCfpxjp07dNcPqchw6t1ED
gy7iiwb2p/leu98jsapMjdIK8BzCaIDpbr9cnI5QbuuTtPpN5mkbFDvMfoxHatTPddikxBwPkZQD
2fX8I8dI11HFzZwxCwAiuQLW31LH5nYZ43LRDRIACjn2d472qVnSKBAjl5aKq1YnFxwGHnepMefr
MVkiiQqwQynccxUndxTfxf2jPGmYLZcKb41XyysqQ989rqJv/Jx1g2PW5QIlL7j99hPG5Vq4Tiwb
NXenmdej9B7ix9CjhMWwN1ISlXMt/zJY6gM/VPWTfq2GpWP/pCdBwqrKIJTocIUlrRhOIjpxzdmJ
nOa0MqnRhupggHixeKtmKS9iOfEg7m/0/cvlDi7SL5a0kEoMM68syX4kagfhzDcUuB3UQXiCGL5T
HOHVNxOJXs9fTD6dZpkHnhtbNSdixBPY73sl4cBEcfPwuBTfeRoSdBu6Gu5w6zgbIH6WWUY4rv6w
txefETmis9QBIB3Eb3RyNf1LjSU8d9kV8UrggQ9vkXsHI7FmGmeoL/Z15CRaaeQw68u1J7cFJInK
qXMahCOPfyE25eJFaX5rTzWu5U9K1JVJ7qCqwUk+2PD4dnETfHr9XDO0cJAkKCDqyHn6HEwq6Bv9
bGUm5UwJrqfqWsUXOKswPSwoOcN1qHoI1dmftVeBslZa7m55/XOvuErDgAUNNtKhxEG4tb2Af4mY
jgN8Y/vscl85FCsT2LUKpQWZ19TYEhaw/taJKbry7CW0xKNpfwiflGl+DZMxC3jIcAaa3HF0mjle
ixAl6YnPyVK4iZlGBVeE+65Tb6qHUYSENCFom8E7ym5fYYGPtbH9dmT8/YiRDRs6ts2sE5diWLP4
u4AN5iF8I6W6xCsIPTlrfzmoHlzGi2QqZONlHPRc7oLkTyjehAvcXnUkggE/cy2q0x2otb3swFF7
U+Jn2lkWxG0/y1VwmnsItJYzXWuXTadZNcLZKflfZn9i66ssQOg+hutDr0KbAy7DMAEyTD6iVsly
VBHvjR/2DwLPDSgen5p/EjYVyyUdw9SQsFF4UJUyrjz52dDCyDO1es5exmST6sKiQnjNI574U143
YM9ji1H1QvUrmSvJXUjgJL0ALCN68vqW04QIXyIq/R2sXlrUA1KM47dCvHHKmnuZtEv8W7VdUZn4
5qCMb1Q0ZXEjy2JeqZyi4NyUr4//fYyEpX43zLNBDYVI2zW1NxgXTMUPzzO3vArR/34+11Dz0JOw
Lz3GI9wDGn/SoAZvu8HRBDPxCbmNPboMFTEeg8diGMbvYSd3lOc6yIT52M7nixgZGvYper82NZqy
zFVM3/xQkHgiQ+lXd9npruDdKR34ovWAOPMk9luD03lk44a98GGR7h45P9MGqBfkBE5so6YZRr1R
IPeycttUtd3yhdiZSRG3X3Wk93AnJeeP08BfkRBa0FrkEVcRGeFp1tWnVYYtuXHkMsh8LOzIfCCi
lQAjt3CjvCnim2+co63FSwiA1r8DNTTx5rsaMbG7jGGknYKgGTz3urkvFkp69wkXR75yJ7h7qfvX
dYFhrTwi5zr5tXO2NNo2ph17IeyjfEJ/y3sR/+PaUjb8hewGPD4bA0SJyLTMWmqGh361fWwecfxq
6JRHJtZNqny1SvVs0N/1jsardST84HIJK4RH5JuHsxy2ZJ2f/hXRCfN/GeHje2NWB7+lEC1nctOi
CWtL5hDO2kQlFdgA9u/fAIUc70B1yCkNjc9WmhC8e93rhy2CBbBMavovLnHaMmKw6ZL7hR2vDwAD
g1MstPsfWcQLvMe5C5oNjPHYV0xRyXIFWWEUW+KUlj06kYKm+7qqDWGoyDN7Fjtw4M38+HklvBTy
tv5YjQPUlOC4BFLdMT4KI0wGnRQXNPbEERAZpFjc7fvxkaZyNF8BBHID6Tx0bITuW9WIOEoMjwMA
Ry6kAXswpW5vnAcO7qLdFo5+EKGXuYIkUN7KAx9SBHZ3iWwtQMyQXLDB4Z/LeQG9fzX96PD+IAeE
QwlrK1Cpfx7vy2rrY0z4RLvIKNh71jKTy3JZclyxy88V1dP/vlVXLuDKdAdj1BdEprogU1vxBEVp
1lTYBiZSoUxjiRxCuMb9dUTXSEA2718gw7ps/J/tPPOpMT+sVigbZImkZ0kJ2eMfWFK93JBkYF3B
rJSPTbs1XEhezvXvIgkgUUsZQRyL35hJVieuli5mxlWvhEtpNwtSTO/dGIiIqmKXaw10nXq/l/6x
+RtgOw3vVHWWg6xFW5/+RsD04PmfCOthIsdlCf7JDKyY1NTxWb0as3mZhN0pz1/d1zD+neOeMKkd
RIpJkI1IE/olIW0R3M53BhSs7cQLCLoITd5UnNOgw1GrrayP1PXF5ERJFxo33agoz2qYKePnclaj
5XPYlQy3dh6HmWsmeEy0pWvMb5lp7eiSRUl8gz0vgPdXMUlNgb+e3vXPB/6Jg44t8EaIZ/cJCJjz
jwfPYMkK4dUVk9oKunf+LKwlVR3fNUvBsPK3ZYgszcKXI8hvGvZTwFlvNGf1t4NeEGGoiOiyn8nC
CGJX5EuhMExk5DssYFQy9ZtHOMDEzbpE3bgp8jCkIubxp357Y3A4QcNWZTCSDVZ5Nh+wXYpDqDho
Lgy1rXqEt2/c24RNVh/yqwER6e2hC1610n6Ln8pmhhM1tlr5TaUfyK2fWabmMErjTZCqv5nLsnKn
qVbNV3WW/eeW5XtqT427IGoX9acYX943V42f7Sp8U0emPu2MAnfM/Jo9aizyZvYuRCr6GaUu1r4P
X3046+igsDxg+/kTcKgkUDDd3haGsL4iICervOb1VfTkPjkmMv40gzjmM3EhUVVEPNNd1pYC4on3
iHkvkvXnjOgSPiz3rwPbnGernUFucR1RiL1FfBb/koYQzumu2c2j7sBxL0lmQu33JygabrmsDgR5
aqAO52f9q+AdP+avYNVuvVTwZwYSVCt2ZnSLjO0rosVgc4xkfF1aHzaLjurlWh3R/Pi/IKdqhzQe
ohVGWKvXCOMgCKT5rInDb1OSxrZU31bcgsYu2tjFeSUngfWW0pz2hZGVAanfyP1RfugMC3EY9Wee
704H1Dea07NuMHuXw1rvs73LrjeZ3FSKTfwfDFJVTf/zeXMWJgkcPQWnpNAp87S2swJTAwVBG/eE
fGQSxdCcp28IY4kPjfqBHgn0l/NyzfCaYFqATpTLrmfT43loc1TlFDhJWk2ksrSyVE27i5gePiFd
fba99R6KuiR0lXggjcN2FiOaUkmv1OVyjvTeOStAzHTlscxSIe8JWE0uuwJgrNVwASgE/HjYW/Ur
25Hd6/y8CV8r2gWy81h4cmv+ByATzfReoNVmeGwMlHTBpHNrjUOK3mwmwjg5TvjP4/glidXZBoXE
hNFNgyo0C/Quee8UMT1+KamlcfbCgfdP4Cm2+KMk9HPLzdBkfDEut0xUrsxl0UgMWk6dtol9xY+T
+4VFD14hoNT6DE6iAn5A9Jox08YZISlPHWqXY5WczRuCzkLpge5RSYurUqLCEmnqubmhwaBnkPBO
aeqoQ8WSX9xVvX5Wo071X2E49NfnT1GpB/ZbGvK4EqAViRVxHk1Xd12B78QFjY9mZ/Rgdv90eo5t
yXgDAVbe/2ywWuWyQryk5Ynp49l6Rm1lxKZ1/ERUqC9QuJkqgoUFyBMu63zK72yU+aHNCOyHW4QI
4GJu8ccsOsUY6aCY+N0U6R5B88oIxE81GerGcCBlvWuiFLz56nq0dnG16ubo+PF/4/ncf3O1ez8I
mxC71TiZQuo5XGgWQIlzkTV7oVUjr+AT5SbXJBkuMKpwNMK3XRSg5SgCTA+QLZqyT6xz6hKNtfyP
bOqCXf614yqu+dDtaDzS2nP2rYM8iMOF+ea6b5fm7Awz4twtVRoaGO4F6KGODp8GQUZDCnl6aXqF
B5fhod3UTFL2c8n5A92AJ/seiy0JZHiLq9u2Orqx/j3gcOATTySdIb7b7+eAm5p3f93P88cPVXDV
l2HxSmiGfeqk+ag6WEBpFUfbSCwZ9P6MPjS69ukDkkrcy6Omj8sjwA1elyx1MgihiWAxPmoicwxV
4EywJRbMGDj3KQNQDZgPNTaekHGzeOuxexW+kWYMi06ExgJiairogvRqmt/vITNpqoTesth8RML3
PcYg7X1Hc691jwJoIN/uH2DxWDSS0Cgv+zziFxJnhZSMx3uCh0myUTdIEZgjyrxQDcHrGZ/cPUTo
NhdcU3oxJyRD0DL5plD+zTfK4Mskn2cbdqxp2wyxzXzjxmElM+ADXo+BBTpBcGY1XPvEQivDQ9TF
HJb3SGQ3llIqHNtG8gkeYOzeHDgfI4gV8XtnclKvMEVGIrH8WMqRcNltxcpbGiyAPNqJKDQCsd6u
q85x36/B7YQK5SE1Dbej1Z2I3V8bruTzdHHiJAgBXKDamrg0C1tZqM0z69iWPVfSVX67a2Luv4In
48YleVc8poYIgSWy7V25eEyGwPeFhqNwjLPlln5P9GOf4KmIUWVnSf/sd2BK+lA6twJB466GsmgD
HxTqX7jJqyguWk63q2QpsBqLZnBSfKSdv+NY+U26YxouIJnOKqdnty6ccwOJPN2ubBD1kqn/kezP
/i6vNVtGvccRgXCurqVd7C1BoBTFD/ekds4W4xmGP2kkBiXq0tnjhIBX9veTAcSst4fhCNf/Zx8f
HxAvi5xwDCoIoRmu053T48OiPicYNGh+qEeBHhomeumcGT6Rus+SSrtu7b1AF7noPu1x018Janyu
D5leQ8Xp5WI8sZehKjpC+1jwlwhlsySoLmBS0Eko/Kolt8r67S1bQX5HJwfmeiZZ3vdEPhLEobDI
rqu85YoucIUXTixn2RN1R7XTH4YJXa+UKlGIIpwCMyJKZ2Cb/jGB/rxubnMybw+yFA+wj4wJ7zvb
W+GLLiy317Msxn6mncbgm/LUQPeTK6qdAkR/Thg6g7yUDitu9U7vXhxMC//u3dTbkdThptMsFVdG
+9gVG0BfSjI87FHBbLMJzmcppI68b612ktD7yTIQB2cZ5ThYQwB+UYdJMhl8QTb7Luhxrdo54oee
B4ppA4If1Tdn4dMvegDwVq0yhhBma64jWZCCuTRC//YGV5+6/KTXhAQ28IYaQAnTyeYo519eg+UT
YX/UhHNF8fewkwaEcXYrxkJ8lrJ5y6jR0vh0mBEbY6fwEieMLwMfr7NLU+4RFyD01xbv/68hj/Ud
owYuQY5K8JbGsjmOpCaBrKT/HqNxagxIuPD5qziGc3ecqFcLlAW7ySImyB/pSZAEbLOK58GFKOAe
5ZZHNtVUW/kJ84V13DcmdxYzQ4t+wMU4UJQOY2TGLop/KG7eD/GyB8UqxqWpdb1sH2jGa5bHySlC
j13MEpcjdZUThgsLQTD+j3Ga2RVPoLYoCqCFJKQfxA7c/zEdQRZm+g0jkFTEy5oiM7U6G6mpOA9J
oS7z6aKdtws623RLC0vPpWlNT7PMjQ9LuI9yNCOZn9nyL1VI8hUrK5szzZB9ox1ds647TZFg+A87
7yZ3FEpr6Je94oWmfYbQoOaZj5MqO0m9wqJiRLSq4/7RjbVM50hsJVZ1AyZUD1r/qLhAIDOfzBxG
KQ/tvpj+REQwcRE5KjwAhmFWNU9AngdZtfUw8LsRs3lQseMHIy3TyaF+tdMvccERIyLwu++0TJ5I
UIGjEqBkOeEDbID+ZccllI1+R2IEU1yvz9lB6AXb38wC0hBLlCv2GJOobnbrTBYCQ/3BAdugcl+W
A2QEebE9MdFc/vXOwwzFPS6T+mjXXVcK2T7IcTL/G/voVLfS2gXc0SSwjP8gD40VPilLcT5IV7za
3Rv7GHBeeN6tS1RimSbqLAg2GJO9/RHt2vflM1NQNsruuUjADMzoRLu6X4NadcEP+ZdPmHZc6pmB
iG4twOVYfE27OGZk7iWExJa7e54abD7mpi4Dx0M1j9zPRqn6dm8MuvKJtMtwePu+5zSXqCnN7UuV
8bLSCYNmCVLBFiKxsFdJp/Z/jVqi1Iuk7Y7iBQWluDxgAhznsFk76sz7act6BhyHUh5Key693VZj
iaLbgCv+5/YyT6LWp+G/NLJQcKKNKJEYdEd7lXF7r4BuPQ21+J9l9PH5eENSNNWtev5qHWm14ru6
05VUE5ke90F0gTPDoxnhQ/1lV/o7iAgj3tLhUtaAi4FWAk8g9ErFly2Fg9p8A3fZWpReZcx3xZow
J41qvaOxF/tI9o1aY4bqUC8K155X1BhcFnDxqBU434BREJ/LPdXMMuFxqgdfSxjcmbfk37p5bYcM
n5qjUQ+dLdxUbSIed3Y0iuiH87tsSreElQ7KScYCPaEPwy9ilhuGltACgr8fMTFn+efUqu4L23Nx
spS20odWGETSu5ZHZmYHoVLNmdm9iLCybzc65+C+XHebPQC3Mq4aV2E2t4eImFIiLZC4kjGnKkd0
wVYGMZjyn7APjXbSlU0tH6qcOmrMqUuqCdu0PSLSHsS2sTQOPCkFsrMhtynG9d/crtCy6xM/GJ9o
yD05Ub37qqWO7FGcIXyrWofvuPbUyNrFghN2x5KemeaNxx52tgzjNOr6Tu5J/Yaj+Pnz8gJxn9A1
gq8H2/PUhLdzZKh63yZ0mR/3vPu5O7B+YfnaXjsAW0oYJBSyVNlBj0FIF+xTO6RTArmZC4Unm0yq
h/CExeuOtpsBNWM/tsxiyDSLPyqQFchpU8zd9uycVaGxv5mpIjU/+ZCteNZ2AgiDnGpDCgD22NzW
dGYPurm4lqJX0eIDmOtNq1u9quERUNSOWG8Bskkj6bkZ3PTxEbLsDgR7gY/l33SB+ANpTMaOv4F3
OpN9d9LwBJ9b8ja01JTksnja0RGWwkBvLauEPzO2t14bpm72fhhhagFk/oq6eyHrPYMxShTbFNVz
4JGMj2gkqf8iGO/DT8vPflVUeqRAh+eJrKMFDhBXy5OxrdfDIrsD4bv8Ai01n+VtZoxBoqwUS6rO
LVN9FN55OeHZKTnaHufCaGjXSTcnwejLHzWDEYpJY7sFy88vmFDjg0xoQx2SsC04/y2/Y0ai7SBD
7OcrhlW4R5lJp2xowqRMaKvK3PbbEg42sqNSSAT6SD660QqV7lJoVevgNJMquHGuvyiTAOvSJtOo
csOoIX2seaMplRu7Tc2NKUtk359om2hB77rv83xQQrdP97SltEtFa6i8BMTH6V4AwJmgDX/5fWWZ
teYDw/pVccNKHRg/AuJMC2o5Qwine6AU2y5f/2Psnt6VxaKlZEfoJ9Rxs2o9lCkKj85bpzruPFND
uMFecdc+w86s4pyPfR23c2OwW3fDT+fYBnfXspakA4V0sLS+4CWl6wAS3cxyTt65S2+NkgaXJ+Ny
s6GGtEbwjl+gb5BsKNx8xsJIUH97g+6vi4Li0v9qWulfyyOqF7M+mr0g+x9osPFatKy4PjnRGItq
xDvacVmfk0d4jrLYDDTgy/a0ojNH6pcuVyqeqyOgLH7wPdLFli9gQIv9hw+w+qyOw27A4vB2SXhT
x9xKDhTSc7vMgUvNUZif4BHqSUtgIhprpXghtqnouiKndhMMwAqm2Vom0Myo+opZDNZqB0tJPzoH
W1qglrHSs1caYNRDShbkzloTuRH0MscH22jmpUNmaVwf9/OHmLj+Cv5Jb8YxljOVHAmeUxjE/ojl
KeHT5SMVJ6E4/Y5jHTETfcm23kOZcBhXMV55/22o1Jeys3t3pRv1LNPPLE1WnI44+JZUrJT+zOas
b3Ox2dUzVZF0jkSPwoG+d8zgGcKmPDITiBKSVsZCFe5sDGCb4i+jShoSmcPJip31YDcXiqNikLWA
ueKt7WAxZ1qp3mio5Oq+nHW5jXc8TdE15umVONxoNybRUreaCCmtJHUGlsC/cF7MXqkCGijScF/x
67sQAJ44X+9QAS7GMUr3Kg+DdQ6Nzj+/UDQRlJVcHvgGBFZy1KUgxLLWHc7N7XPhQ8wil0Mt6bLd
LqC7JVhsax6lXKZRaDYzEYH6I5lOTMoV+4dTywpQrsI0U2PQuGI9YVrRmbJPLZD/u7ILZ0T/xbsW
phPC7Di/56kloj4ajTCeayovYruloCuXSJR3hYw4kcttUxhwcLPvJImhHQIP2/1WMtzJJuOFYYGX
Oe0iU/yc937AZgtbSu/e4fEHBJXZP9qJKg8zoly2miy+wlthtFy7ECIcEUrbjrPDSfRvkoOP9O22
Z2gVUNPGVpPJyuAL7ocz8mFwxIqo9G/ZVqHo+tOy7GDF75jFu8fNmvKijJHPc5mCQ+nDWFlDQc2b
ZPIydePHacRdeeA2anDhPqANHMRMQ4+Fu5fyE7yKoF8eZPDvRQMgfSQGX9Yr9g3qRxhol9ky8e/N
b+NyelPt/3QosU6aqoQ/8dF+vBl8RM9b1pnsBUqEChpIPXMyk3jV3x/haNcIDZehoXGtz/1XJfAh
guHKOTsAdxgTIOLg1Nth7LkOeLcKAc+JUMVkJtG49GNaSrZfvyrLO0m2H/KVeot5V+5F8kxW03oJ
23CTxTnA68bpaX6E4rqDAndRsek2ALB+6huZRQm3Olr3HJS1aBSoGfr8ekqo7ZE80/K9UjeXahff
GJjKINCVHs+vragerRyAPsD6y7HtacgsA5QRS7hzoJzrEsf7piFySgyvJLIcgSr9qpf2MYRauwWZ
+U094LdUNwk+FdrGscOT2Mj6oidc9K0mY1rXekujF9Kk0T1ukasoZflX+JjpizE83geSr9b4xtin
SDxcoCZf/Du3GmVlXe+P2l/HZp04F4uStSCtrf1h2RkaRx7l6kscs983OgMIk/oRJYpQSCC/Cxvw
b9yKW4TZDS62Mk/zRCOK91+BcSC5Q5pYZuwzEUKgLBd+DxFG9tGZCAo4sxg9ljKFlUKx8R3a8BbQ
/l1OwcfjoB+hVhuNJ90sYWPrZ/i+bPhjBmbiOOG9u2A9i8Oi+TE4qTvqKf9/QyXMlYebACtBQros
OCl4UnExbtvJYsTD/I6T2idZWzk1tsWJtXtgsk9RkeiVW4/bqp1HGw+wP5pJ2w3W4SzOiQ0AVXUU
5hpdVvkB3udTHVf/IGAJ6ThhYsekY3kn2vcjdRirAoTzlQ6JjntHuuTtY1E345fZc2Fbw5Log1cS
un24NrYqKkNFc9sayb01qQpDe81NO/1QcBgDqqAk5ZKNSm1TcDE0QaXcvUP/N/Pu1G13LXSyACN3
9yDInuZtGsIODRyHr4DcrI6RnCK0j1vSoBAXNGXm24bBus3eh9/0RDQ2X62Q9qfDcjhDFhXg8NOX
pbBpgqZIVHO1d/eTP0TTtTTY4xktHqeB69xgg1KPYOrYqKZaGsSWroOUDNmTw7P9l5H8++tFvYXx
TUv0xYxKlxdzkgSSQ9qfHbKy3hGGiClqj/sDVJD1dbV1B1YKhzaGLuTnJfHDxKF2gAUHHjvKZs0J
RIqLQk+UN7WY9mCk68rGH6LahpEFgZ+gEEMLl97v3DA/PyYSCkzBH8RQCcnUbh+376Vfsdo5FRgj
Qz5OCMS7CzJhexYKHHLc2fRIQpKRJKIqEt6Za/+FmC9/yVRvX6b0n+t9Xib4USxNuftEKS9HdqGa
/Elh9aJdwfHTWgRq5HUePnG5KcaeJ9peFkEnBKj1fWgJmpX3zCZDZEMbIU8bA3jSr6CcVQn7TKKV
bpTm1xEy7ynF1DV9ahZMHCXa7NNAlELR4iZuFPS0bu6G7cb2wsNzLzlGUSubiNCE1F2lwQyX3lqV
dVsUObnZDzxFH4xMN64uzAZ/482GHJXESk6LZD8Vx9cUt1glOaQlhpHqFLTXLE342pUXW6ejlgZ5
hv4zEhvol6URsXfBemksqstO7am/ASfAo04lJb7lalpWqtx7dFzlHRn2bhf2gCsMg5EzLVV06vHB
yjpUUeR1YHVyDqCGS3H9X6H3Zw04KOU4CMpnuolMxYbu8ONNM9DZcrsS+ahFPjr41E3dNtEO3/Ks
mt/RFX/IymOp0h1V/QokNuwOJA1vIAlyrD5NtamXBBntNZQDeNpdeyYriH8ukP63WGagN/1YgsZ2
mfdZB1jFpOMA8vdBWCngP1ObCZukX/69Ll+ilArW5PSk/rGGcXDkdiZUrvH+Ntfg02Ya7elPK1rh
oFO+ILGQFcv2OHnjWZDmfy3NU0PH9EpjVTL1F8VF3R9hCLOgFrFL8BGrxO4xR8BvLJeqgI8in/rD
2h1mMugaYNRElD76M7dxXdD5IvIs5lFi1115sxkp/z8q4SU4eNH9AYODG2T5D8thw4ueCa3l9icC
6nPJlLlzzKQfb2gUdahDWdMUECP/S75c4RVL43ayC1hTfIDszwKKbHgV7Lh4GfesFtHhKqW2Z5lD
Lg9ToDfOqF99/O1cJpJuIbqnnkLYJJH95IpAnwr96t19zjsOtAETtvfhfKsvD8DYoLc/kHNdNdRy
4W20BhcV3XRhy48fcKCYgp7nHSxbQmuqbP3UZiBbt/qefmZmw4JZiRqBT6xIYRpoHCdNsDJ/nBIJ
AAi99fiRXntaooLfGwQKiY6HsOx3pADqtmUSRXF41rUJzZFDsR73OEFuq/euA+lsRco/zOzYH8Zv
Rj53aKJZ/9ylW1IQZr/DjNCguNpJTd6AndQJHeUf3XvLZv8peGDqVemPwm22WIW15sbfI+Dg3nbl
3lcj9G6bb5h4bKUG8YmcNR1gR9+lj9xzYxa+enzE70vdFZyS8rwUrFFgi/EdZf/zP9UqjTgR62HA
m1Y9TdGnPm/lapesHr7u8kh5Wm+D6OQ9O7bdN9YGIi3CUQMUtNy/8AhKvt1BKd/H1/G3YwpFqmDC
V6b1GGxAtbxSsMeHGrUWpYwot/bYIZhszHubYKX3fAc/n9oB5wrS8Ctb4DqQNoQ4ZyqV7uRGWOTz
rSlPAyWzZQU+0D40hgesNQiZChXDgZIOX9zACapBribiCFguSZn0KgvdjFOI347kh2lIC960Zd3v
paY8e1dH/1LA22OBP6biR0dPahuwZjwa8mjmPqBvuSMACGrs1SHzC2GVvNFr9BU45bM3oZTyNx8y
MVOhBo8puZJj5vXEtATyZvs3ID6HYnRXmtCgYtdRRDVZZ7Vms1XaNGNN2P/2ykNutbzfEckZIfZd
45EzZkV8wc35NmnirrCpfcUmjQbZeXW//bLRSfxC22id8W2stHKFLhr8Qdoex2SpKlm7OTwnq1FW
SHSeBHBs073glgNCkLVto6Mm8va9a2/kTrKJFXty352X/MUPo267DwveqssM4trnGZMDZsLa7A0N
BlKTU0QQ6d92zDrm4E5QN2T7oRz9Y+O04OpWAyzp2+BzsJhi2+1NFWReDJ5773iqdg90rQZ78HSL
Ic5Po1HNm9dYX6bdg8KbVFWRrMILthK+CnUPiWR/eeGn1NY1PR9vp/QtvjJU9rRdxj44eSmUE4l9
rIkU0NRogp8hqsGZXOoAO32XxfPxiGCOhgiJdU1y1gRCETYiC3hD/Je8xf88kRkc22/x8EXI9TYD
GcWSF74yT/qh/TMpTcL0R5NnioYn8sZKwQkQJbxHdqghBOwBsvOpFEFJKkTNddLIzJ0wL581X1lL
whwxwixJOHPoh72Em6mz+k+ORZ3H4+tAf2FpwaJAXF+wSwCfAlEs4A0cdlq6Ux4aKxyiobcQtjy7
m2uOHuOXR3N0C5HGix2/S7q43CC+fB/l6iWp53yyjN8qaeIGEm8tX4AqQCZ2ke0/oWEgxYPOKX5+
fylk12P8xRWG30D4/KYX4MPAl8NHIaxJZuFC9T5Ai8iriXFhz+JWU1oENEDMOpnpGut9kOuo4U+A
glgsB9q+mzAkpW4DJ/787/IcuIp0vgtuRlRkTJUPY24ksQJuaLn/IHmYJPHKcL8GBzXe7dli1IPw
0LcwddEzm24o5PAxwY6I14ozGE4qj9+6Y5XAoqYhN8zZuh6eQW1znm1uBIBxjRtA74bwTUytXS2x
Xj5tKWmqNMHqaEBFziIBcu9AYCWbxLjwpxHkrUc4i1FUw+ZeEUVpz3ery6IRisIuH3nzSJpkrOn5
rnEIhi41A14SBr/ydie1MuJrMhtaKe4P+/VGjTTXU1ME10UvjGKK8kEatHtVgBExuXoJNKAqFDBh
IthKvL474ul39TeyfQuclkAYIGPPQKX5+y0ffdUIRLXc/oXyvj7073nGlVTWHf4QhGJOvVHHWfaC
FiY0DYhrAUzE1ESZu9laqCuzwTSxNgQVHhJvU6CVVOmvTzAvqxQKPHtucd0iLR6l3HwsAOhT8JjE
RBtcfPT91mi6i8g1saotxILjHFnZuOEQFA2oEwV5G909GbiFvhFBHrDAon37cr69JPuuJ2HYiVTv
T3nwFrEmFnKzKM8moJvKHIYq3ZfnFXhrrlOUoa4wLkWYT7ATMyuFT2eblQ1MpcVc7YQRf/lP3K7R
Wvp0nTN+L94subxPyiZOKiB7RULSY48TDzUz1sjaZIiijGTXi2CAKfDt+CnPF5VqVCkZg9aX0+YU
yGdDyXX98MP2L7UAH8y0lVt6tPPXgU3dGrVUmWrWhsIUmnJA1WhsutIH3S+mWNYcxDj4nGD2SueY
vilNXfPN8HvMKG/6N2qUsTPMMfQKW1VCqve7yUZUxrgowPt1YwMzcom/ctvOlWERqHstL+2XZirv
p+SH6N6QCh8NCzdkgR7+CnarWr8NkxTX6Ud3KdE3zwCwKUxFae0ob8uY9QcN71aJeCE3SNu5Kbts
zfDZwG5ZbPDRekWr5L2F3FVkf8p+i9m1pMIlfaIW4157W5AYL2TOH6sGRRvf1kFx8UKh3kxxGkjn
2g/FK3JOIRfQCzOqtYUNUKYKicYRsuCa+pKHMIgiQlYsAjOuI9nobI2n6lG7ai+OsUBpcy3mM+rQ
322KwQiUFnoPmaIcxghQPx4liFIznpLfiCXAldjun18ekuqs0UnhW2DAzS1J6xViIFQzvf444FCT
JIo13ilm4DExQ3WTPpNgkfqE8WMdGVkM+znr3ZwQafWi9V9D79dmTZxywX0QAvG/z2FAhMoEFPbu
Eh4h01hGE8MIuW8o8d8YC1OYcCNWsSdeKqt7dzgIsU2UbjJxxmPxS3FNXThqAsm5R7sBt9hdgzt6
Qi46rNnP5wnuF0u7UZ8yA/Ez6lwlhZImQxa7gSOG5aiTkj4WS6SmglF2tstSZF/s5f2NAI3A6Hz6
iA5JnipGLRmlzZoxX36q0jZrnM9Wy/jFl8hNjNSFtveeI3pYXYtF+TUiW9aW7pfej0OWXPV25Gxl
n5K3Uzq/yKCIyOpbhuGFre+202q/9UK6XE9QjlQA6FOcuW8ukc2uWwdx9m9xom11Z2cnulO7H4jO
Ouw9ssfsLd0ouTaXlf4DHE4/BT49TTrSP0HD1WBrhaGa4XS5LxdqJ2Q4HpHBXxFIJrLkLG6O4znM
PbCTbjlIP75kW9TPStKzxpAdRosB9gDC1frASJ8bewfu9sTud3IB5IpWbK18ntYG5MIKLJNuuBLa
k0NP/vf/IN6py16RISwxlW3CRvjv58tgX7UzC91wiEFzCI/SQ3wgfpFLHLIbZKJLyJr6UquVlVDS
h4ZAhurkwY/JQHYoWW5oXBtRCJCwXfpvhAxb9pVzvpDd+LLGDqerxGP0dJtOfcuOp2ATfUb+wffx
Ld738l/3G/oecApcrQqc1JQ+ej8WQFJNCdnJmtG3wQz7/yCns7pMSeCv+lC18p8r1GkdIZQCjp1G
qFs/L7wWyiwhVyMTXTuWfbHEZJ5F1ISO/dlakMhpHirYMJIepy4TiOvYP3+fK9RAfYsg5RaZugak
602pxopCuroX/ZrL5pxb6hZKHttg7b0pWSQ0JDNIQALqvL08yl4THaoigX209qDKd7MGIyMCUPMI
Uvlp0vW3xwk47lnY/Pwe4HMnHj42sraeRe5PBmdgQOjjl3u6NWH1RMB+rmqd3GD/xqrusDTcpXAe
L4dk9cAuJ7uIiT1Xqjj8KO3tMT+BjbmmgEyjKUoEVfiDuSGPvVLywwSIFyqeEgKSDGNESiFoG3PL
IyrCj1ovqfF+Lf+m7QhgYfRRFymzy7kOtg2hf0ZuPhrL7lyt+qh/ghYqQ2Fn4uNYQayUPrADi+3r
NtJbfmGjwgi9HoXXfyms0VqbAQL/dgvsYCsK6ZaLI/fy0ovtynGLEMCa2+Tv7asj/Aw8hWHggSqY
bdmZ+rRIKBSDbkmykLiDr1di4oCusa8BsF1l6pVa0g9qKEoSrd8ligK2xMr5lCyTEULo/M7c+c8S
Ip7BzCHn93LNrJqETus5NRyjjy9qr2PCoAEphokLqg91Vh98408WUsl8j6ygWyNPHGveqH2eCaHi
wMGaaYqKOk1PLSTMjDdOkXfcEw6Ojpdg8B6pfErjvBICJUau1rDLAPxVhS26SSa4lQm6zwMuabNc
pcahDlIdrtMTlxIPlrJXB2XUEvwCc5gaP+mQq49BGqVNR7Vzkut89sOvNIOnPfPqeKaXetuj3Pbh
23ZxTHfHtjG7Zr9mMl0FsHyse+/hbsg+ClqfKhrMvEkBp5cNDmASsG7SoA3BwQi2PrHFRNb+LtuK
Es5WZcwuxKEU02mz3jKMA89YdhIAvmRzWZEvb8yd1Nhw7cCEEmd9MOn/ZISQDTDk0f28mrXVsCwV
WFgRmc+EJUBWUtjhHxHmJ8NukKxde2jaAbG0qJ8FuoX06UDFU2rYkVd59HfdUifIDRqwYpOXTtPK
QoaHOWsxodQ+Loay2nQH46/y3ywB64DsTAZY+RRlC4bt11Jl7wDL6wietQVQsktL6hY29ZMqUu7s
7eXjwslvZpVFX6ULbHLDJl4NMXRgE54ZOlsLVjf1OEqZQbpEa1NGekKWz8YGFwFaAxs5/Gz/D01a
w+yTTY9SPv+QUX26d3BeCPSaCHVIoxIiPJRb7ggFFLDzA/yHeY0lNxs7o8i2+uLApdqDglD8wbr5
rRBj0IBhYreCuDpN+uU/5DLW42PdBkpWEz1QqmthHUm8PgEbLg/qPyiBHyA8q1CWUNTpu4uugHEF
vOqKNKMcpQe7OT03Ck7fR7Q4nfIBdQg68KUDCAjhw0rK/1NeL3QN/noEtQlZWl4UWCn+0iQh6KW3
B3rcvJeKEh4G+c51kRidKGjq6e8NzClMzcFncd1aTQyrShQBDufiUFWLbe63tKL0q7gesuKcXTDv
VFd8Kg+r8wqa1N9Aagt79mm5Ov6sIIV/Jx7tosmbJc4fxbCsFZBau/4vhVz/37n/g8bM0Scqn5Jw
dPpT9sFQ+Q6cJlcd0/MYq3AZF9Miskz5Cn24jDRWq93MtvgRFDSldKUyVFBePVtNKjfpS7ygiX0u
a4gvE2mQoiIWQqWgvgBMUhb5R6qEKfK5zgutgDUvZoQ8ZayTIqOS7smLrA9SLa8ggc3/DtmEHDYp
0zpRT7dWPHvq6XFhPLPYado1es5lay6tdeD9ZwSZkvA3mM6hquCXqlpwzdaWaoXar4YySNFPOA61
NA9AhnST7RTbkN9OhoCsgnGeL2PCDQk6O45IRX3PwkAjaS/VWHYfI7cXyKBqU91a4nsfYsdBm/C0
iYyiPMyteXFNL+4tUuqVwUAm/PISLqZdjHU/Dtg9Sh78ywCZj7Xulr+SxooU8i8N397VTuA+LXrQ
rGYCjww8+G3ZYk2iKU5T0E3ZFYFyYKie42TM3ebX3fOr+0w7FIrBpfLIkmiStV/W9W2WPrl2m23N
nyVat+MRBU1b24VDutED24qfNv35oXdnOJ32AFuzY0qOcUC6W0JjyKg8kBV2xK7BP2Rfaw7o/UjQ
Zjc6Wkw29f3itV87+i3HCIV9uwdEVYDANY/j/xGYYPFfVOKdcMUDKahxveo5gHil/CdTDNmDKzuN
1cj+R3bniwuX+AFD5VWSXH1QvUYe5SQGm51uWmcsLVyQaylsUa1oaN4KF2JXP3gsJROcq1U14Clo
yiTQZMpn16MO4bIuCdZN8oAVofsnjbL21bZx/Ft5ztLqf2xsnG6R9bX0djXJK7vMnnTqYBnaGkyV
S+qf8oJ2SomxpgH5FVA0cBcBuyULBcq3m0jonwtnUbT/SIsuuTBC11YhLQB352jixrqTNgeyhlfx
bj0OBhrsg31FP/t1zUmUZPLkH98k/uzSUsG8bLgfYIuIbin54hQQF12Eu08r3EXkhfD/183ubgL9
P8F1R9n1VgMgACqwlC8CBO20YYK9/lgVTq4R1gpD1rhB3m42vMaOw7HZKZf+GT1O4OkUChj8+0nf
epgXABGnDzrY5VENGUkP+WGglr5nxHUvQBJMJHocChLdrFII5WcZ3oN37Mj8ZsRyYw/Of3ZinVKq
HTPt2CkzvghylR4g9C0yMXEPXk4wEnDGIfgRBIfYJpIKK+qDLjDdVBKdOgBmfLZisjpe1qWwM2PF
JEGBITTV2IVASDfA++U5eGkTscxQ2iT6/Ji5SurYiCpD/GGHBQ7rLRvU9Fny1Cr/yDgzgMx9uI/l
5DrI6AqidwrOFD3F7iZeg9RaCITWndWFNU41i5/DyVO5j31xhLxBkIHc56o1dDqhtbUKoC/dnwg5
Jxp5wkxUYK4cnG11bxYFxPBl/LG2uvokyJUJ+OTx8tFRjNf5L5LDGoPLSJyIgOmfKyBjkRc/n0dT
1YB9JezS1qYTLJHaU24ngw5mfq9lQRpZ8eE+7FhEGdEbDBIpq3311fO3eUq3hRhXRk/pk6Qt+CmZ
gzQv1muI4/NHikRnHiEYGzgyInZ1kySLjvgRNW/XQsIQUL9bxcpy6NeGhdLjcIuTk4PiatNi52Eh
ldwAgdxF6ot+G0RkwWRtjSoqboU/g1Bc5zX7pOo+yxTNpRD97fxuk528llMNwwYKuBgC7ycqKPY6
qra7XTet4KcHNIrpLwtYoolCq+eeNsYOyQ0KTwxjiYfyPfd/rMdpTnaWYY8Kgd1ch1FHpJeb8aj0
w1SnOrC5jyaGK9y+WrlWi3v9nFjd6ZV6BWMVK5gp2pn2b48X8T/Md2gCdurxbbIXLiizAOXakUf2
u41UsIvZjaV8LNBgPrSaeQobDQful8anzeRD5z80E2HUBlpQsiUntPtQPCb4dcS/+yV+ILRrhc52
IpzZFiIRhMTdJ1RIPaR5wKGwEnjKVfj31LU2V0ylt1AM5RSq1LapZq86x/6kLCitttHqYtUtPpNi
R+wxzM4oAEb0dZXxJ5M+MTVHyrWjbsksM+EWX8ltB/E8O5L6EjXrmX7/RKNTntBKIbmDHK/H8koS
WwX7CiNQhN/j7TwTmI7h5U1geJ05SRi8cctnw9Eno87S1tODyJWO2bImmQ1qLeEYvzq+pDDmS+eb
h3N0VSxO6FE1iurrvT8jYoyFVrUlevF0UK8sPWFI14SWfRjFN8CLMBsm6YnBDH4EupBvxDpIHfvJ
Ht2NFGaDgp7wheU7L8D9bdu3aBBUZjK8UVkFCACZgF75Pi7j4oTxpfYIyTcGOB4mKopgyd0SV//r
V5FtkjZrIxYenJkZYFcKgcXZ7t/QxV7pCBGd0U95xtLGV5NWX3eUy5zII6x3AusZcWdi95gKo29V
JnAvwxdEGYw+EdWJFr30si6BEKO2c20sso7JQS8nf5kjjc9fBqF3wP/SQMOwChKc+jIgndp9a8aC
gVjalQAdz1LnyYJ15wDftwpOIrKJudNXc51TDX5YjmMSpL+IlCnBg9jG0Mv64Zf4NlKSSCWtPbFJ
eODWdilITJ6vKwyoQ5NpgeJDunx1PUjHpT8gaPQspLB3MUaHiDi78PDgsXqVA6Z2ZMk2aex1bIOI
miMghNo1LOQXLvZIYaPHQUMYuOrCa/7ZLfz3Ujgg0e06yELdqMMx+CcAuQqLyzAcwHB24T77jE1L
NozbKa8rGmq1BVfupc86/e0FwrdCbFL7yozg5guccDtUd63xB0veJ5OTaPVMeyskTEW+HIiVhCuN
VP5qrecVmT+LtZ1h+OCJaPEcVixv+G5TvvKkoakWefjMu+4/fzCtvJVwFwpYG6BCJSnyz1VxOxow
X17+0yO6oG6KNwfwt0bMa7xmZfOTB416PQPMZL/BlY0PcY3rw7jFrNjN6rzQvll7yfKIdE59C+EH
1kAF0TFs7BpUf0SxLYTVGCglnq3jcSghNePPTl4Jz0mT82gntyWP9P/QSVlWcAlRmV6MH88jX04J
emDgUIaUIilLBOXGyUxwwXv3H80aRTE+sQN09jiIrEChkNemf7qd0ZzBKbpzd760hXF3d8eNlTSb
15R8hL6ME7BObWpeabRSU8v2wVHyEKGLk65NFVYXT5/LXfxgvjQpkE6oP07bEj6mAv6PsK/lxzHn
DuH6IJejVJpDNJeJJ5nCRtz0meEr3IgpxTSnhp8Jg3Od4qA4SDYfUvnjCZubVeTbQBtoZNGsxjLy
KBV1TX4dZ6ulag6D79uKpjQDipFCwsfLs1xlYpy4AXFb2B+pjBnWb1FD0Lfn/6GFHnFcW/Hw6sMd
K44agQOtCobPzo+vrfAweDSfoQ5C44TjJLI7xOLoaIFd5VskOhk6rYAGvBiYCyBPOmIc/d1OM/D0
80Wu0tjDrqVLZWAGOM44G7Qdc2Jqxv1jhtgRyCVlnQS6jmhi1FTbP0JAE4PS4dpWp758LBpIww7X
2/lb61m9oXgipT+RWdvPevi36LE6qAFuDfgzDvWMNx/KSDE8X2uzYlw1a584usDydnXGUAkUUzXh
lSbUmQUEYFNOG+d7I3euqwhpNADuQbt0ic7MTlmF6QBLqnf/optQHcT4zuDuqiZ6wigg3sll59yj
XXam7LM08ggNhE5JAGL6PEqC3Dob4jVhG6fAtOWse45siaDDaziVrmdT36F7iT8a6VrqJRu4PxY7
+NxHyEni1w1nbcbVH2P00y8UJnUEhV/llTN9hG3TihzWsu0vCJipcJd+krX2fN4nMWf6BpKxcToc
N46+31qVtZURMANgw8vbVjdXPvxLbGcxOy9t2q4C/MWiI+mt4ueUs/zTEMg3INjJb3ADopknjZyt
pmqnq2zhQp6sMaFWo4B+Z50M393sjIIa77F1NRLY9SGXnZQLp2zxjrxi7LT1ITXOnguB9HeEfuzZ
8Mq9N45yzbw6lt0fVrCcC9mD75g0lqvN2VoJ9huojPBMgIcmWSfo+ZR/DXdPkQUnmNVG4dzCcYtb
6Ea7prfryWYdpj5B9jnOaRgLzA+zDhhl7QlCOcXtsvRtDxg7WYHQaMA5TOKPDo4eydEczXsUeoiT
H8pybHcF3QZl7ft3PqrIKa++mLfxP20IMjm7zHb0/xxzlUdrklIOSUylJ/wajjR1uKf9g3bOcPj1
Fpi1427GpDShPnYHs67oHW1Ub0zJdoijOIw0DGUwsR40ViuJ0mruiItkhFbJVI5o0FX9D4wVWArc
GKEl2/uc4NiPdW8FRIptTC76DA1LydDr9HbpGzpUrKjGg8rPCzlbDUzz+zKZFoqfxKBbNxHDFsc/
r4j/Z/U0qNoiZtZaiHHYgfwwGS/Obqy8Il6t63LiZZVpoRGxflxAEENOp8uFXexsdR5eCPGnrZbz
ETzbKEEhwaYAG7JDm3vVCxF/n7sOQiy49haPjXegkM9w5GrPlZgMNXq4IDa+BT94+AOg2q2F/BtN
OEXIGTF8QMxFMq+F8Ck/Fc9XBILuQw1mEkSahWI8Ijd7JxfO4qv262EiNaA2rznG2eL+cMxBssjF
Op0iEvlH7yQkk871TcVzTtPJIBcD+5sEH7v5JRG3ajOtyF2sz6c6cpufj6m30+pLCcRpF9CNDFIq
a5Rt2+aetcU9UFtkssqZV9Y0glpwv0JXY6iVcziyeXHn6vLPFcr21U+loecrtsAId/LJei1NJQD5
YnK2OPX4evaQNejYEyuEAVeVsPxUmc2DTXb7vvwSpiRZoVnablkZNvWKdlKii7C2qvY949jmf3vJ
+ctrNgmA08qMfO+oCoLm4jrjyM5dhMGtHjlCHLmURH0isKBw3FcBdZOn+lmL5rWk5KwBCtENnKD3
2tKXPaAeDEsc3dHj4jkRMX7GZZzU+fAVrGG1wL8aZstWuKtiXRkXstfPrxUhFFXdaOAqZmdUiyWr
23eJvM5LRabRjyVzyNTEnv89zH5wvgwBQotmDi1xDP0U8QQFzXN3QecaNw0s1LctGa2B6Kjbk+/G
uCSNtGJkQv9yw/MfPnu5+vkeIp9vvIX7IWjCtKToOTo4dC3CpM675cItl4Jv3gdELBINLGxS4pvn
oiw9UfsJoH5UMx//K9+yVjopkJMbVDbn6mopeOJvWcvwlT9+Vx04WChFHB6h+8HGl1OkJJp2P+Qv
Bz5wcfIGaIwy7kwoXNGZBQIIcVyM3GYWk4/Nu7xzp3qDMFYLn9TqTSq3udN4NoROZw/ECA0dUXf1
Ss9/hvPNTmhqR5eNSGp10aXa0EdfH93WKSTw7zrjaEvzC8qMtrwkL/FZezIJeAc0CaLAV1AbyLPF
0NaG8YG7LK9so9pRvdVlUFMLOfaDOusI1+oGjZmglJG1m4gwF7zSpWQtjP44pN/ly+aeB7ndmF4U
b/r9x/efqGsqyfcw5CB5CYjD/Q2tlsT6UlUcrHmNOYFmF/1qPBRovpq2L7hBJqSyLKuPp4DVlgnx
2tvhsy4hUWw8dD6A1bptd1AByYTZwf8YIQ+5iz8FH8fAipb8T+gj/fv/yDgh5h0awYdSEKhn0Trk
KntCTAJybDcRByI0nmI+bJ+V54UnIK9mubc1NpnSL1/ot7/6iKmzNBTufPeLoNytAmFU41tVG1BZ
erH9nzhNQB+OveA9CR2Gox53DN5JF+FlVjnXBW29ben9vDdENxDnJX7UwFslX55uWOz/T0s3dthb
bUg3+v89qQ0YwRbOLcwdwDzTQhPRaK+z+rDLDMjNNi8SJzJGNTjnNNU+eNQuy3Hhuu53n2kBwBN6
j3OxOWAjz80n3RPPsUNTSd5JX0HLRWa0k6Aq973G0Unhdf1iknx4t68iu1LTqGDUZ9Teq/ZoorCr
PR3lEMXu/hHNsk7R8sQ8dBbs5pAzsNudvoXXePX8GdHu/7gAlGeD4uYSrz5UV3gQmIIxGKTHKrAi
J3fazF6b0yvOvu4fNmVnLFZnxbgB6blT3Grk6jtTU/v1k1jE5w0gNEw1rZZs/78tLnC5U1I0fDnv
wzfeAyCJPJxlJQSVhFivtYDuJVh6uzUezU7A9IZqH2ouxitZEwNo3y39Az6r2oOXgvVaqmPy9RDN
FBz5YiCWhe/NCHn8ZIskEIpPgAHRwQxIbYKphByw7Z3xj6w9HlgmjHMuIc/Yi4tS0nBIuCyKDp3G
KkaIGAMsApF7FnUI/pA+ORqYC/uNn66PA49pGxr9a2VcGweAgxUBcRVGxVsFqr5VZGpw4+k9oclp
Ec/8pqHvkYseuMEacpEdRkabsLboby7X53ZxFCzsOPU2rY0DFPmcXDaosED5eMIQCoZJbutu7QSt
Rlx3UpfFLHe9oT/ICbF5PyWG5Whb2ujVmJLExIrXljTq5j+rdJc0tG+Xy/gxGLgCuAMvkS0kUlQy
Zu2RuAathxbr1J8ivsOuZu8dxa0F9+PhjmWvEKYBbhc7S6N6aGaLK9JLB57pNkziqZSnGB8J+Z+N
stQvzXZ/GejOXOMyuFwZP1oPSAbVyphRCbPbMZHNG1UMnO0NPTSqTVrEKbGH+TkiQQ+9S58zQIqo
b7tahAIyZPr55eHV746kkd1rdokynF/W3QXFc4WpR+pz2CJ1QcHmHabC0BlP8C57JQNx3wiRRoQZ
BwptYhz905hCy+qGMZFJBUwLbTADXjx4uPm/2HIghQHYikcncJp1Iti1Li91hZRCaPpkPX3TM3qq
/ipXP2Tk7tTPmVfr+1mFV7ATlKG8sFdwkXi+LxJgW5z1j0b9mySrRri4dAnniYZilihiEgm1dcnn
2Z814JOPGBbo5YSVyO9AXv2id7PgayB/0P6F1hrn7ygUMUtzoxK5d6+XJGqy2GBDEo43xZ+p8r+b
SssDvW03KV+YYyXn8iZkqawvnnn8PYco8qsbDh3aE0XY532pmSlzs01muyy27mBo11ft6vRWgEHo
Ivt7eFpH7vfWvzU52P69/rTuudRIG69ZpwbEWIiTlwJIIYAZf9+Sj/bmcxhAB6KjYoaJzKRrCxdq
GYga4bC1P5orebC7nNRa4MfUKoae3eoRSKjanKz5gymucaUhEy0tDl7tN95aowR04n9UtaRzHiLy
lBtSDnDFAYlhiXlyfzkSr8bHLa448GbnqqJSGH7nNmRTGyHy6kTfrfj8p0mB+uVLn8DKIhjxui+t
/AsSiu5dvEMpiAlm3PZBfSlAo6pXmdc8jF4r+C4ZqA9+H8pH71/0CtomjvgbHpRRpb683ZZ9iur8
q9+HoMx5ZqjBInwNiDFZldGUFwh9wXnK4GPAYD6ZcEutqf/vf4OzkPhIqMud0XXvSrzxQFisGz3Q
8r23IfInwnwnE21LNk+rdXRi1NUXk5ZniS6tEWCEceWiKWaIdhiESnik/qBzSq42efpmWp+zaldO
11Fb5xNe8h/1BSQGaZh8Myxm1zvM0+uxcx3izsWJdbNI69+ktVCKgFb7hHuWoorNQSwQb4s10zHt
XaEvFT0sikcOZIA5TPDyuUTiZUdueA92pL01zlBvlGEuqSwh9jT6Ez9qip4U6qC0H8gV3DC8oicB
Z+R50QEIKM5C+fZ3q9xXxEcE0UCidaRXg+Z/m3L4+8+p0UBikuOrqzIW884lbXQ2XqPRuntqRff3
CCxLrFrpYgRZH7Fed+K52GW1KXY7zQns8Vuc4XVrb18J6IMBnWlF8XDrMziRrSxPpJQFipUxFDRM
ZD6tIT1FzJjydgl8cCtiQSL6ea8ZWAZP7k1bF2NNNksucl8EkXKQm+jsT4IpdpbPESQyIloXAdwN
LBpvs6OqPj67Vs4jFjEcGcndCBoWk8TtF7spmx5IMrk5LapxVMPiXTPBVDcIC6R3VAWg8s4eYazA
8codB1G8VF4CpkZ0DulokEhlociuAfSaOexmGocRGAgTX+WXepz2NkxooHXLbYCexx+0NJAOq0IT
bDV+IP0UZxbVYr0G9E0+y5pZKOh3v7m4PjsVLutdXrq6Is9WMAS9Ke7h4Dkuo3cITIPo3KEyK0mR
zt5ZUJUgw19vHFVlsQombN309IASMncUYC5CsZxKHbQ27qTkQPI4kM52MTgfNJIPMaL3vmbW5IHf
KJ+tQzyLUa59ge81S6ovRdXEpd4QEkS6NQFayoMkSEa6y2MtRHzrHYyk0VfqkL7wH+JRj9CdUDKg
X2Y3rVlGiCWt5g+Jtr8isaCHxbQZmKPiz5tcHiwN+9QqY0HkUWJnSa9dqmnkflWemniSW+vZBA00
KoF5+X6zm6lRzkHVhdjVF0JBYngZAW1jZj3AkHP2ZeLBlMHKT4HfxrttYQfnSu+SeV3sAmiVhdxC
NNkYPQ8HZ6OXMs5it4P2PU0SCi6LHvSoZlrEvVsLBtIIdAsK0jJpXlK35IOAQrdQ7fJ9D3VO+r4p
yT1e/vbHRyXrbL8GTNQwEI8cwNusOZCaH6WKTYleyj1FAwjI0ZVtKJfnVr/W3w8+fb9zpNpp2Vg/
E+yPkLaY3mbZzz+P2XXlVgc5B+A/sjmYzcgaZrxAV9awYkTdFb8esVgSDmnbaLLniI3U4v8rEace
UDOjtCAje5YRAiC4C+H5fSi45TKRvXJQIX52dw7biuB6Wll2gj+Fv8rX51i5Bx+zdcJZHGHtFQtW
hYsPMQ2r47XgNXsiN86BTx+NZ4iDcdsqE/0jvkRKOkzzNWZ0DGRTAcucDKJdiVYz29vujEKkqRCc
vSpIjGv/aZdpHzFj9O5KaiXRu0Vu2eBP+BySHrS/nJCgpdT2lrnomIoZVj0BR4SHyuCThCbkvgoC
bTlfoyIKSO4dtw9LqNv/AJLa1pzgMWpDuKh4+TyzkhTRuIIKRvxWKY7758mDZ8wfmg9cyJY/CGGT
IgsKVnqSOXwt+RaSfFcqCNno18NVi+JLJLsnOcGL7KwjtrsBJMGrljhr+atQp4h/E3yg4WhTZuOm
HvHDfZBqk2i3KQOh1BNb0Ov94t2fWYVMiWN5VfGdxyz8I3nMgWoIOnnen8T9QB0L5RfOb5dYQNNG
AigFUbgfZQ8mJ+oZmkg5z3LE+QZj1pyTzESkAUH2ZrgpBwLOtIwMLhw5dUMXXcuvTayLKHbkcTPq
bAQlJzbqjt4c4wqUHWyOX8Fx0toarku1cwfUG6Aml//mEOmMkTKQVdK5veEE+ty+92hH4oai2GjA
1rmq7y67369u59/7Nq4qBV7Ub/Pz52M/t0GrbH1l9NbqHESGnzhF8JOI4nAYOoRe4FaulCv/CKMH
I6R6G/7UwEW7jziB5eyPnczle0EeS9+/lok3djmyZh+ooZtzGv4GVMOiY1vR5hBtT3hMZWYyxXAg
K/J9KpQYdn4YV3Gq3y7sdSzrz/KYx9n3W9SjmkilQOnwC2T1jN9e75TC52I/Wjscdaxt17M3rs/S
yAfCY0wvHXu3vAxWYzJVlVKx1YSbrfDC6M1WmlYQQQqDHHcSw3yBiUAJTUYiBSz3zk0Idp5T6iOd
19mF527mW5+AzxhwFidiYsn2Dsa+Wx2UolmlQTsVrkxq1Qa/5YfzFvAk7TdQ4HwJB9M52sg9rHn1
GA3rpAN29kcbZs35i1pcxSJKdfZgJyziNJQPhZbTbCHtXm5nsOCPyv5TRMfCW6LvK7AvgHr4bEbg
oYiE6VUJckyAZFgFhKk4jD/Y1DFJ/vzhL0l4iCRhBSMvA9qzgh861Fi3jlGDGCkXwOdQL+AsD58U
BTyUylYVLIT+REqRMd9I0xO/zFvxYnxF1bpnTs5j/9trr15IRTj4wTu+BWI4v4DxPXaw5KNaDYiB
h0Nl3V2PLKafrLygQz360ayp9BbUfrsd0dMduCIfBh30CWX/Fb7Zc9JMMmFiXfCjQx3m/W1i7OKT
rDKtXPkICAIHbmjkBwCv6wh8OzuEH94hFH1IANO+sptKMCVMs4cLdoy9SapDQIa00fHCXh+XbzVv
ngEyqEkWIYq2VRFHc8Y6DsnjN9CessF8U/C8SqlguC6xSgzCLz+7sUajktJ9cle4vzp2ipX1UKI8
YvMKj2uUTNjvMt97rn1keHcaVjIvGvj5VjSowRRDjIJPKUP4+htzKU3N2O8ZfVZOux4nBtVz4n4p
VeMEoZN5cU11W5hE0O5kPYsDKqELlY6bf60rQBamtfUtiEHTn1bMwrh+MMot6eaVCPIWVQJuZslo
YxnrvGgY3v1FwTtzalXClo16XF0q2yu15jrDmyUztxQJZnhGH699exWNGveICzRwOWtN7Iew7c6R
xPGIqroWn+W2K8654AIBGfIAR7ApEkqnrNQerJc4DNZRJ82HPmCJeq0HI6r3mhqIG757YXHASv5i
PhzZF1HBKUHoDgF2mX/VFvFAGHCS2Vk4XAESHy/+rLx3qMXORMDpL9+0g8DIScrCKJFJ7eHc50bN
rE9ZoFhCoTjLX7iy8Mr9BzTA49TYqt78r8IGROEcwdvBxZDWL6UWi/d6D7McDSR29euHu/vmfOqQ
MLbLneaSrGv7t2qj6wEWxOq7kWOGwRIH6pyiNGIX7jUNJWdA2a6W5CwbHCOL91lux7F0T34HgDu9
wWV/sp9vlEC8n+RGFgfjAAepaUBMdLfq+I2VhHPdLUi6fChNFqA3DjuvEWi7mFyiOIxH9DOxm+SS
a7td84COxByMj92RQJhPLNnvi67nOrO8AlNWs+t4NuswBluSHPgIpK9unG/ZgesVc3KfD6QKTa2p
XhByWz2pD93WZf8H+cG00X1TTA8cGXSMgGTMqFVu6d+CVDOW2abJi1MxhM969kfAal1Iydy4Gh9k
UsDZcKphRB+dT3y+nLVLN214q56PyKvZ35RcPjS4/sZvJQIrRtb9NIzNPyo1qZN4OTCdQ3mZQR2q
wW44QGe/XoSSrBbF46daHuDb/3G/pDxjPO1uZGlotcqUHr8GjvMWIbK1E6IUgcIRI6Qh5cmoxXrM
i8BwderHk3o7a/redpVH2y1wqNf75G79uV+BqMg3QdVlJb9tHNiCvw41VB/rvwHJmeM0baszcdR4
yM6Yao1TayfzUHeBe/ShGmJ3Rb8Kdd6XWgnid1VuAvkrCOL7L5X+VMq9Yw1SJjg3RFSUy3ZXLY2A
2wKfm3DUmRyI4NevWB3LeXjGyPIO6DTMciAn7OuDdZkb0xiFD4zMazbYVAPK3Kep/OJDYZ6lX71C
j+Cz5zd95Dh4NzRPEbbbcpzYIT0JBLFeWYBvU4OQkhl+j6MBwPYs7mZ8AokvBfDwXhpp3KOKTlPz
z8mjMV5RrFUBDJfkSR2V3Evw3e3n7jgecpTxsX3uvRhlayvzY02Inv1R8rQyKZd56F62L5XCwDce
tvd0W6X7pBOcuM0fSAxeQNU0xJWsUMD9pJRXRkBbsJPTRuKBDgYAL/KZT7Wb5JKmmwsQgYnyzhC0
BgRxHKxlAw9DO5OZPUh2/E1ynufumD22cz9/HU4+oK5u7r2CyAFBLKIMBJDkUApJsx5GEVqSKqQr
DkBC2eqsuoGBbRMOqbQmy69uZtsuosgX1n80brLvm7kvrzAV0FboGFR2O2UcqpwCgM7jwoXM6I6l
pVdHgkGFk+seV/VkGsdyavb4vdvZH40D/fcT0h2X67LVOkzSIBDpDIkPAqj9uPLR95J4qu2wZ6F6
jgXYwx5lA0AIWjCTBSZ9A6kp1vl0l+WjAIrBkBE3T57A1+hDL9FTKz/rYOH6w+J055mxeMxzSnI4
olyeOcv7/Vmeay6rIfY6xNfWqKnNm/9JV20ZVmB2Q1ZREn8BVY8uyo9A/qmIA0GM46T6HyAyf6Ra
g2U+vxM6agqM/CLoaofEKanUqq2YG7iGWLdXzLMemWz5qlmON7JHvJhLy120QhJIUzFxg4Paogfu
C/iV01jFq2eiKovh9egF4ZeDzxwysCEmM10H2dWhIMMc+UPqGlv87GUPkUmITlX8g6d6ntJFYmZA
tKReXqW3C9zFsYZBb2xdQ+orKDbtLgZbj+jzzefOnfJkkw+SDzRVai5vSKm/jBWIOq+5dGG1xgLx
wYh8WSBeiNAugxZ24zJqu3xgDDXlAsWjBT78pmrTWPRHMJWEK05ItRd9nZWW8pMbZgai/bqE/L3m
ypjNxlrFmKQn+Sgs8MoMipMCotDt8D7ZS4MwS0jI9gEV2wp49geryVom3723ECdaq5G57ihaawUJ
+pVA4NZQnWOD4QoWJ+ZX5vDiKveBNbdRks752GJIWTboAihC4olXqUQqXNDb0LWNilJeon5aLQqJ
+KkWvwQggrmdqVfJgUQjYD1FpJKrxAUpzdaR8j64fyFTjhglmWhtjFayFSuuXlRjAAD2+UAZkAqs
feLocw17nuFSWfkKgnS9HOZdrXFu1IOBDsuUp88qp7GoTDwjQLIteC4FNBfeZm925HoNlwYUuo7X
XwCRQDAYXdLfbaSVf3g83bMD4cFlNYtAk3SMVK4Y/olQaOf4AixEYYXunQfTavQ87RvDCjS8TRpQ
CmuK7ttMPTSBWBy+ijx0gYQ4mDeuThtHxgDT5Lpuga1/vG1WZucLLf81TzKFm6rPWCB6qZQsX6jG
IY5lZ+gx4feWec8d9m+qTGjMlhEb26PHv+o4KxpqvtBjva/eMe3bQFXYkBRBHDOC782XO2dpcAgg
EoKbnULS0IGbazhfXhFoH0qiNFkDa9ndjYJ22dLuKIQxJTu1USnxcQgUc5PQbCxediHH3NPpFxSf
vnOcExcEuY7XIx5j/502bxFAAfohc+v9GhDx+zKtxf1mn/Ak0hSpqNAXEx63VYDp7zzFA2iUpl3x
K9Bz9SsoQKc3xxiLlyCHPSeLBLmOrCFkLEZPF+ZzMP3cOw+NsOBr3BrW+P1TutithMsVvkFvT4K9
fxgx+cvidy9OcD4Rzi3S2xfrWEbIe/nEUNIPCPiGA0I434u23Vz4B+JQJS3N1N5vhOZjWE7ugLHj
y9CnLnajhZzDKTDO3HptwfTY6SoegQKiyiuCSBRODZ3732O8y7xd4uS5ouO373DLcpE0XO+ISqBs
NZrRXC10uGjqgksdij+COQSbFRytHYwO/ElWMVR+NFvFfxWVh4YCyixClwOmgfbBJ3kLb31B7Kkk
lx2Oezs6i4Ftj4+q1KN27p9gtK++FLYJ0UMcOPkuIZYqmjbVw3fqz4A1bcjPH0QHrpNLdkqr6Stn
sjuqd6/6+9yhqmVAOl/2uOHOtYCM4LeAHojLugI9pZ10WOKzcfS11hda6aUMCfAUbBMJqVVO9OSA
O05tGMsXpM5p+E+rDlPU1KYLsdrUPB53LFw6moXqd7Hebs91cyuhZCHjJy9PNNbcFn3fgHK1UH+9
QwUJ0lSQkaqqOr+XaUH1mD/BUAfLfAD08CLfiZGQCpksVMmUvIcCyuS9ArrvXwptvZUgD79/h0GD
uXSAyJ6wdu/zNex6q4qsG/oH9iV+VTLNbRjvAgsimJ+jQcNZCNjbU4lk80IVR1ytzXvGRmXefpTN
0Eyiw74d9HlixZUHrYgqdM/J6qerEnUJ64F55RuPq5biGZPMcG9dty1lCI0dp4u9zDKvFrW6kUau
WTJ28QhJyiYo4UkWzFLgqftRsJfu9ogZcgHZs0wbtj8l8jT1QaDKokNR/3RZ+zY+rUt8vLhgViBJ
P9fCGLDfW5OeUl03eL8STiWwyHiC2Z2uCAHXaqpgHTUR5H29Jdiz1VRD8Gi38qF9ynJZuUCUB6oF
8TMmLC+Gb9MhEWHZtbsPlhpYHlGM8jEdGcabAcf35EqNGuI6TpYUTt7aTGfrsdsC5RdZTMew4jjB
1DqOQRHHVvZOAoAKS7pQ5iKntPqXplHHsF23UM/fuI+03xRbtQsWQguz635SoKVDK6xjCzlvnCVt
Q4LQ+vg+v1Fq0rcvEV9QeMffsNaquCt6dAMi/gdH3RWagKhJPMl4ISAANEQXDYLsWXsYbc0LrgcJ
niGhQKVE+hn/gk9y/EPGhVi32C0jVH2ViSH3kRQlf0IodugwqtA9nId3WnlsA2S4repQ2oax5xtK
I3TyPFBR0yTIFoGaOi+ZUy4u0n6iWA5argaQ5AcE555jOgbUuYmEnoCFl91frGGQAOBIccgK74SV
DAKIw+NTwXcn5amHsN1T3PN1rFU5pSc1BXBGbhq5DuNzcaXgVD7R3RygFnC0S9/DrJf3rU0vVJ0n
H979HXUQM+c7SugEmqk1Ad7mQjck7vAbf+Pl3OjQnjzc4aXvzCegC74hd2QTE9I0FTsHD9i3+kQQ
JtCmxv1doMQOr+AqNRF7XKYK+S5m/O9mgJ7OGZhQkVM5FQpCT/5R2zhxP0LeKDxAB2awybaDJ5UW
jxRsKF21pGWKAPFIJRqBlCx0mMduTq0xcVXh4x/X3ocN0OaABXMkbD9NZLDrrU0KLAjRXKuYHbur
+CTyuTAHSpFsCAJToLrAcFizz5nEVvgTdJLLFw3/5PpcSA3zArFGbVpWf5/y1TLP6YoEiyvLOBe/
MiKDR24V1fXpknIaaI4mqTbe9iKcYHv/adsiSsz5f6Mpo6ZJDF4t15DTADfhLkyLchkLDGYN7GxS
1XzdPFpVJZhSb7ndax99cn9iWcrPnMsy99KYWR8SFO+gg6Ae5VMPtKlSvDeB0qESfYKc/3IGjEt+
B8FfFnRFfBtPGjiLO+lVmDdz+F0R0SxBTvL6kDtUOsLhWNQm4CI/bCd6ifJdtc+lwdUBx6QbKUXV
KpJaQf13KaL8WkjhWggixRGjRWmW1VwJnSvc6OMVCbvwLJUtWHK8oPx/vZMbq6x1qMfemy6Jzq0V
xLrlnpAkhrhvaAw8/vZhOquUOI2x3hgM/Zl9Xb7cyuhexVpDEfg3blBitryXfwsNLaJDoAK4HfaF
cq2axIXoXb1yWH/YGAUHt8+N0eSrAqfVjrqWJf4NaY8kRVUhMSyPKaXsFVDAmB+i1KQMRC+H9XJt
P+BU+l1I+1dgMVKFq+GfXj/mZfE1jqT3wtpnygm88rf5EWt9OZlx6xRC7ndZekkFxpCxDspguRAp
jSIP9Gew+XyVKaRiMiyMCPiBlvHwqHoIs5bLuvl74rCqFZU1SflJns7UlOdujmxSmEx/hrlnx/5L
vfyGqYAitaWs7ipeKV5QhP+ML5EetecD4lsBL+48dqF7kzy9aUU2yM8UysYwl0qdKULedrVWhC6v
qo+NpvpsbQYo+Jm5kNw3YUxiIlFA1vCzkdn3c7z1wY52GgjllRhrAASqwhWKYZhkr6hxkmwe1kn1
r2IfcEN9xE8NmenYFV1PXUgwo03XZPXPbyQwrVzQBiKeFdagP/JEEKnMz6FFdFp4304F4pUWTVyA
kE4G7kGP56AdZft6BON8Hb104MIc28JglG4u6osVPxVccY3DyqBvQZDfTw8hAPuTDqs8j83p1R/c
xZrkpMGBknmVkAMTHkPFk2yln2NHHk8TYWTLQV76sfZ1PUxq9G4IXAPNGh0zjZV63q0OarkloPSI
chfu+RCdWlsMm9so/70A+dRmz1lVKObgmjCsUsGOZ3yD0+/rOJRoITyMNm1T2i6/2xeN4W177Ftj
KBvcnmd8BgwmHA2TywxRUnucJGuNVLBpUpSDyR0/TYcgTWKQwKF+7ZRfibIS0mqebMf1mVLuZv52
X7qb6b0el5sXO1R3G3fWIxJJm1FHpRHNvaF6tRbv8YKdpnB/8j6YuLQlmoDPXSzVybOkARSOjLPI
L/sZzFXZf0l7ZRbnY0Vl6m7o7FsNjbZsR6zdnsEWTj4CM8y4On0uvv/XJI+LMhaKFNit4t/d4Z4Q
M9rDa/v0elgCLUZFv9hiRhx+H36WIYQH34pJZ7hX7upzPhYxD7tEVhJAxGtJ904Pyun1Hka0hgLW
9W4SaiwRVBUqPelT7X/T7vmbGw8UWO96Tpo/yL1MkBZyyetu24EhbBYS2WMF5zFgFQ39g3pBPzFD
okI7A4YxpjttetavoS6ru4RAORnKdiwkLI/+aj0hz4PyWvHTFkySXKrp48vXmSjQUTbnJJrLBsd0
R8wzXY4NgnNPKS6+n/1fbjrF8drgeAMFddIMgBa9EGh+7cAdry1yQvRYrc8ofVSPI9W761eUOiRW
ncILZiNtXBlvelD6Bm6OooSLYWRvtKJQwiW+KnG4jShftnhvA6YmUWX4iuIlRN3euIu2W4wOui7Z
pw1j+W4iSw+qeOku74RfaEV7QOveow19R1+3xMQ57+sVPOFfg2BoVa4ePEEtbZQN8W/9AIPQS3eC
vObUe92RP7qk//UClWUvCQRQisWYtv6eEI2dVBw3d+drcglO1lKmaxn/YSWejV4dMI+SrM0VDPS7
3D6l3+XdIQL9nEs5MrtqQEKIF8mAKFZcXIR6SaLkRaI6fZuEWU7kI1oPUmJfEQ3y55N89sOM4b5Q
pH5EhaTso1dqK14+AaCjDXDfjB9Re6Y1lzppmhQ95LF7xUpQAoE1psfXQE8PyQun74mGRbWv+pvZ
82zLY2uWeTOy+OgqeukSAHME2dsBT5WSQUoMTd8e6kBcs/DJJ12791jLp1EXa+XjFIU7+l/Fumuj
+YcrQZpH+yPsaRlVLxqMrRt6XTBun2vq1I1FY0ZowSRTqkx3O5pyM46npdaV7nuypw+SKGsKzfx2
sREyiW9x0blgdD6vq7TVesZR9HHc+NbVtRRtppvmJ3Ezz+kfJHTHKhrHV+53hDDGQJtDa50hIinX
018Ha8uvKRNHh0k95hnhZUu8mfpP5KNNLGGNav560x6X+RJdVaDiKwygfjV6619y/wB7Oo+7D9QM
yGGAxI+ukcXNY1aoPhCO2JfB68+XCGxmdXxK1Rct4JCGT8AOxJ7bvjLbtBWqoiOwlWwJVZTf8yZD
XyaP//RDb5wOARbYunmL0X5bG+2d4pON/LmrD0e2uaKinB3rsXX9B0DluWkDni56FLmoNDizP9ls
fr7E/ucP2uOsTP3AIXv7zU1HMOrPi8dJQMFksJJK6/cxFPC9Blc8j/LRbBoIcrnBv2qDcirgtTkf
8NRNJw1D4vAB/xvuLNdgR5uJ84FmZBlgRvMqjBCjiXV+4r72LMmr1fzHRFaTj6Kz0MbBWh3M0JwB
3a/Y0pV/UcDs4N7lhB0QzvNrKRnik9cy6zE/HBCy8sdk2Nlfvc4ptVMVFbKIXNFDMIc9Zrj6QoVM
UIty3nxm8ci8c07Effjl85mklU/NzLCQvaI0DzowlQ3gQICwW+z+0pZuvNNd1C+bTF9LUBY+clnF
R/Z7UXVnNAfZd7Gab+1czg6dw/kTch/lsdYOaM03sNojcOLQQRChnLyC9BtZn04WEnenFjRQduis
W+h7WdLGjPtHQxxWRHtwm9usJVF17hrnwUlbM2C9TsSFb9UFKUkEz+REBSBwRugaNwN6NtZnaPMw
EiQzQfjqACB337y6HCgkp2+cn0wK+OcH6wOBeOeqty+L4q8lnxjUV95muQSyb8iS8r5G5IyrOIi+
XA9N8kWBHsiSkAEp2G1Nyb0s8wambg12o68fEc/vhZK8z8tL8XpeNyj22eDO7f2ZG3cWtgELKhWm
IBpVraNg54YfcItfOiX3tLHevPpeON7XekQIcYs7fh7KKKBEsAYJPHEhIAnvCPOhkTJ+VdFXX4TT
n8Uq9ucARhprF8eLtEZWlKQ3J9gD8VSQMfyVZrbpSiWTnp/ft/9RNGCVBY91n+QClceRRZBu7ptt
/iv5O157724No3/bTD93ARwdquMChmwtzvgNemwVeEqmeNglT+l3jUBZx9a+UynIpaXhn0qyo3EB
Nsf/Iu5IP6CVkB9/x+jZGhXL68IT8cxjQ/u3h5IF7SAFXPT1jlbUzFx0u4RgYZIYjIIE7P8pTC/U
nyPVnqj+Du+/DFJI5hi0tW0NDwPFejD0k3uzWUz5XqxjHihjK/hbtwcHPtWwiijAn5nKi3RUwQnK
PUdsFDmXE2Pi5GEHBq4WUdtR+6RVAS16si01KiFV5zlNuUKJDiW+ImsTIl2RGsP42+rCPCdh0dkU
2wuZwES/kC03H6rNXEz0Dw7OWr4ONZS/6SRoVbdoAfsBF+T1Qn3MmI8FVzzP9zeHunYZ4Mph+ila
pdjZ70+jxIIeiO6HJgbZbGUi8dNse5yK3Ejgr7SN/I2BrvRDfJJy/wbaQByoCEjsEGpNM0hQkCbv
6VzyIWXaBtbAH+AM1QNtCJEtjhpvGDIq0/HPb1CnpHtX/cHheKcEUx0jfVzATCKCW1nWfU0FLaPy
LX5pRyAvcG8FNJnHNZ/lFpjhe+8D8zzK1lAo4ZIye7U0LCc6s9SYEd6o1Q7yUJve/Ky88Bw9/Ox4
kIvPqm4pUs/LSPY8vNIHdQYZD6XcPV1MPpTNz0hrZesmDDZdD+ddrSDjm8XskyUVbCAjhBsp09sY
UgNFD7rI+B22Nf0PL8Iytz67fyIkPg7bPjEKqcaQ28KLCHPSq31851KSJ2vXYBzvbq+t8P0DO383
DuYQrdVdTmpC+XGXcFtDwhsVfXtiv4mMf8snaqPzzeD/Wq6Wc3avuBaWK79iIQE/9Vi31O6gVY8F
9Lr4xL+12aXwmc40qRDYz6NKGUStkwJa+dmkG3cKpnHOIwwXYI/ibVjWKXWaZ2ARG9TSDTZCDmnE
CiVnyk8BVjCtW+rLYOGlsJu5sCx8cdNslIdL210jHf3MoEK5KWdkLrQr4PINbvafq1hDG8wRSw3i
MQPn1FwzD2y64aBqLrep5fjqWAGmHmUX4qIETPbHdOyRxbe3u4ooijIWTKvSOVkV8ZlHkRklgqjO
FmJ2M4UOHaQaW0FC06zU4OnxSEWvpVvdZ5TgqROHLwlWr7du0jYCacUXmsEToB2H8YVJkEGD/qpk
eAYEhnXXLMJ6qG0qaAfHfmFjvaZWN8K6TJipLWOB2imycIkcjv/6Wz2c6wfEAzTQCes+MTBllhqv
GEirVdR8eeiF1/I6mgnybtJQafmqd23iCP1xXSIZJ4reqwyL4QSvL5CNroJkhEaG8FMCcSliGndu
wptc60jS0ri0alZM0EtSDoSYwUB8rGU8DN2ilF8xDkDFE3azXEVAZTLxegm9mgc4ovb7sKdxAhxW
Jy9jCmbRMxKpxTLGqELvNujcZxjiQEe4Ko/23N91SndLgRaMi9fLO8/HDr44yyDXbawVf55IKkhs
I2y7RdCzOt+FBUxsIjxqynuWO9sECPOc7Evhg049ErfVMdz5hwFpNRfjfn69v8ogIQfDFPNEhWxO
WQkrsVYeboOSTmOZ86bSIXIEt41ygaDdoYoIL1l/2hp6YS5lZiRa2EUWxlSOLLuQ/DeeP7kS+wKV
T4wLZpfX/o9y6auEq/izRwyXh77jrLPMPMVf1IXBIeqbM5NAkmXAzoylHrvpG693Dq95tJF18T28
S69/GUBRaxSeoG8EQOAXpb2yvjzpqYhZs9yyvOZmKX+XUG0BKfHMe4AWjE+LnU+j0H5Wk3MQ6WzI
QLmTuOtXKbRsowK3L7gKtCfcEyUg/Ho+qXN7qIPkgu77Y5ChVxFXjOzwfZjiD2ldMNW1nULb0PcW
1DaXSbFy4ocsF9a4QEfl6xOZqK+yxif828k3FL7yZvt2iMzAllM3N8HIW0Wqw2A+mBb+1Z3FJ1IX
QTYMHdHkY3x3RbXApu0RKGMd3WV2f2MAYTquEPIxR08S2jShfwl+Au6jPI6SkAsEg1q1Fgm/qyXD
ZEQmPbBboY5OtJAwkMlMmiNEFCFM7rKtbGb0YLMKCWxgtn+5LTxE+azlj829z3/bbnv87eyllYb+
x6CEnjvXrXlV+sMZHWeIePVwFxWcTo/JMYmTrQV8qP/hOwieDRqUjqtYgeHx06YqdOSohVuLTlW3
PR0P2+KazuxYZZV/eKaPODuNwzYxGLtOE5q1ImezRaA86+gYmyw9rrJPl4tUxsPnPUrwpGRD0ka5
LtlZLIlrYh0DJ6rUM30GLqQqr2+cbuBJRb5xMiizLcLXVZTUIRFjaItFjUfumxj3KD2ED75s83yE
9gUn3n6bunYI9cPUAgBDCiuILtJfVQqTh//n5lyHqVTGT3Ph2pG3xLYD11k6zXpdMa0iw6EvZKEK
gOL4Mnqip/vsZHOurwFpyw1jSw1H4o5ziDd4qTiGlBPuDHDa6BzSZwhwotXZDkM2pEVjaquQCCPR
U6mzSKi0LTu2wPfqCC82QKdhJS6s6cKWfcM3FNyhr7Pmt4/+ayNuw/rP+eMSNJD0l3HONnV6L/St
ScBXqS4y/DemXH00R+tOE5UkGdJwvy8rG9y10/JV0FLIbXlb1k4OMMTtgFel1VShYm2XvyUVTTZL
mjSiFC8jsaTSz2kvbzWkBdtRTYC6hlmlwiTVfih8KKE36OV1/DW/to2MTLyT+WVr0ogihpkMl3QI
2f3hwxDqE+iQvueFDdswxBNwua2+6O97D/k5tct2hJYIQ7s3c3rnP52+oRwcjuVtRRDZUPmoNs5+
3eJXM3RTygt9Gq0x0weIfRpU1RYs03P7lO3Aq5ylWJ/Ia5vM8bgSVCBPsov73lYNpH50CHqkYo4+
3f55kCzUPHRw/YFFlCiBmn3olpsZL2ocZ7y/h3Bb9pExbCEXev8eoD4XssTnfBGqsvSSqKhtRSeO
VMJYyfiZ9O67chSYaiL/CiDA7jtt7mj6dhUBgDLRvkiNDzWZ7HSdUuqXtmii8Yu1fFksKhrfMCge
kB1S6k4ve1NcHs1amuuxJbamOFcg/NjJLW9ZSfA/JXOOoMYkRWPwXrM2ullLkv5w2L9jx5478tYY
VtGIvySFyvFkNv7UKOxLq1s5GKHmlj6pJCjmJXRWSGPRgd7A9t2sDgle74Zu7eeYXSqtKLZkNqgH
bvcfOQ6uy2sgmCeWlW9351h3KlJ023DlcP08AsrtUrVQse0Z/YKsw1vSrPMC/XGtbdR2qVTaa03n
339PGwJVrMAXNwgnbr60G/cEI1X/989Oc8bjb32xcdnnDQTnpCJ6JEhW3YTedCywZmzau1zLL4sk
bHUoZzje2r6t+23EHN/M4crmR3611R8thYeYlcccMRbA6ggKxVvk4TRiu3Ubgim0p6LWEtQQfXSk
mK63RqZ3n1gpSsC5K8Y2cy+ERyRliHxWlL/dFbdxcdKhesFWdPPFgCKH3aKiNf4h2lfrjK7yNMp1
EP1SsrFkVIZ4s+MCnv/hw17c4EOEWSlOOfWG+Be6n5timWN1fQUgaLV9QrC+wUkdkrp0UbnX2cXG
E1pLOS2nRRy5PEqdA5GsliodEX3W/VWqAtNeJEKSeeJsMmmYfi3bnvoxBXt4J4V4ggKalS4nc4he
ZOUSsWXL/lTxTOqv7QZOr78YtR5rBQLhrCy0RSVs1tRHcgPWRjgTgs4IoEznzflStstv9g7RyZeh
Z3uOqaTnz7TXLtnOC8wKcNzhCEidYB6poCbktkDro9hPpmuXhF55iqRtpto7M8iqdi4rdfzZan2O
gOiGzXTMXHq2m7amBHb9/1rEaOjZTRomyexwxxdld7fdYzRYJHhOxMDZhsi+MjXIC0eZfTnjSw7r
EITCD9+WNLtvgYs8sWYM9ua5SpG17avoV1498uduxNKP78RXdM1C6jzniFpo7MGEF9a7GP9i3zK0
pIkhSs/KbQsYgJLeTPaAXcvTg2ctyB5RMe4EMI6Gkzcv5oO4vYLMX2w4Yp+IvIAAlYxx6g2hMyP9
NPWj8ayNziIZgZs3xcZSra1L1BaiBxLFyYPkFfmkLCXtUnXWHsdBmY3UDMorVJ+QbKUzm+pF7hyV
O9xIkz78i3+75iY4Mm8yRhUwV47DQNrouN+Zy4qjoY/mG2RdA5HHm0sguAxbGaI5ftXXFmqotULU
dIx2ITth3LN7BgH42vLUY9EMPVwen5iZ1+Y3OQcLcJPL4U9qfY+EOdhJv+ymoFnxBU7XPMyKJNdo
RWxe0IGPED0h1dShPf2aEpyu7YRkWo3HBOZuPnVgKnSf7OZAQeuuBwmk09nJDaBwVkSsOz68DVDY
M/rpasxsqZuo7oXSaiJBxA5gmS7GZajPq/k44NCHczrQpJ+ugWIMIyOErAhc7pT8JBY36cSt0CdX
CZM3MFJmacygF2xOJw1V7nBWqlStR+MNSD48uVCuzEtz3l4jC6FL2Y9GwSnYxo2NyyDMCV4QG7ZZ
BkBFtgKuF4mC8VEg6mm3vbI9tP3dBpiT8+6s1aqC0zlP0JYYYk2uWJ2e5FWmUZqdPGjjHc1KkzKM
bR2aMLo7enCQ1lK4truZWlMls14giEoKYVuI9hQwBdH4lBN3XwFA7lMkmg21F4zo2mMz6KABBLru
JnSVn4PzTxyzcE5c0PfWOGFvyrLk/j+BB++WZFv6huK+xUE4oph8z8/lrAqDalPd5ZMV3HAbU8Y3
j4lOm5qvKn+QG8Len0XXkPJ3Q7PP52X2/8XjRqAyJUxNnxxrqVZ4dSWszKlq+2RbC1v1eEnR2MBo
9M0b4OQ4PiPQq4/lUBh3eSOgzhU1dv/6Ge/VnawqTtYv3ZqR7kT0FQ1zLRYnPXa2tHRApO3ENt7p
yIK9UMMX66jh2F2M12XjOD825VyEl9Y47nyGUm5hJ1CSzSr6BTlE4MF92yRUT930thlJGxqLDFwl
FFfF1RTLdOlZUIjaF0EZFbnN2hAOSmO9bRsuc4XTlV7WORWys1b9SX6aOuhzzTbjEk8NugtMzsJj
tTckCds2dBOTdToXw425X2smryJZU/wGAiMh2fUJ579N/flE/GDRzyOeQgBgYm268t5nMeh5DrT3
jOdHAUMW2PR4vEODp5ndMCQbUubfjWkpp3vDCLqZYCWwnZkFjXmM4B3tYTY4trfwxY+CmC3mKfmA
hq8WEcBSXeVtNZgVavTBpWTizN9VtWM6wygRkLFoE9BktNAvNnvzKgKiSriiCaPtTkFM0Y7xYTOH
mChRW5geRcCIQ2vOIrn68oMESV9m+hTPOA654I5vVh+vtGuL37TWtMMRu09ZtQre9R3ZLvOih1eK
OUgAtTZk8+HFb5v+6IYAiIQsw5ZRj5iSq6joUrRjIRH8Jnxg9JsNtyqhaBhSJHMljasvpP02kRUi
kuZOmQYKGbTyY/lBfHuug0jFGosq5WGgETRg9wMQxbeUId65Jml7zHRGgDnYsArfNhtuOju1Nu6J
J90jsR3NhIBmKhJLkZN8/YGexSt3Z48pYahZ5hxZpuGQdRPwXDNe0NVyy25xGV5Y8FpTGXAU7DqZ
t3ZljlAVTGaawJg/p5zPpPjlI7IuzlwA/VES0eHLu30viKB6XiN9H7zSQDuEOc/by8iYrX41Bmfb
pDupLJYkmIlpb1qPfxrtpO1laCmPu0/4vd4lwfCSoBh8c2S8u3kJWKsz08R1myrqTeZKT9Q7O2sl
/vmxWs1VxMlF/9mztxu7Vd/z4xuJ+GXPNaHQq3crLfMxcTkogQoLLD1OUuvicJYFKnV1iN9M4Xjb
1cxDFYcznZp2264oiWI26+RL8ZC9eEvRJiVOEeWgnbDSUapNnXC3WNfuvhxHAFF1Gk69nSPnfsU0
SHZiLd0qaogDS2lwbU9ImgXuGsbC7MvVv7XMarYC0PF7v9aeXtofq04JENyErYo4kY2zWGhbAibE
bb1PO0z7wNaBYGVzkpu0jr9JuxCqKI0sldh2TRYnIqsKXhPEYCVTcTbnVB1DjdaHqjRSCCS0l7Ql
Gf0QATrOIMXTF85vc3g2PPjBTQdqR6WpKjv8b353vDDpYOxDXfm6uiddfO46DHtJILd95sl3jpjJ
cPrvWdNu+kw3wDJ8RAZLseQqsoK5fLgBz0K46H7JNXRLP6s1Fvl9rIITDcI8dJ0mXwc3dIvBLlge
mplxPTE4TxReG/S6VdO0PK0bqcWyyZ9rIuY11FjhV4fMIk0EuWsnNSPwJt/Qbml75//ulKYUJnfv
OvK3zvVqNNByQOSfVw1KWpBEH5ngzZdUsRnaGS4Z4tmjfwaUy+bKgd9C096EgJaSOYBNCWWwx2Y4
oh4seK9iAVkxCj1zyANrs50+Ct75J8fAHUcLTCX2U+YH1S50LdADdz424ZrOUL+fOpkBz4rL0F/4
K0rjmPBfnajyd2uhA4QSt6X7PR9wfpNCmZvHGHzYIAlponzA92FX1O6SzBVfQTNM4onzSG9KeahF
4j9akhNDJEpSqlok9zG7KKqKVgytCeRqcSIBqSNIbUde13C4AW6E9lfoUzILSK/h7Nere97cSeN3
DwOuzTT9/Fr8sqcYHoL8ZZ0IqvinmTrbFHeVjgY6PhGanRJ0Rgd9kwtMQuaneIKBAYqz9HHK7lSs
q9rD6d26cvJwgH8I5OloXR/lXzZiiy2jq2aNtgtzldY6CeDei+290gf25azvypjfVi+GD7wBDW79
VEA09lkzSubQSRfXhaBPtk1cLK6ajN8A9LzMjn8Nd9CILLCzO9sSJRvkOB/FO6EclLdXn1X0xIPK
WaDzyDECbBWQ5801pRCj7L38A0CfTXxPza40XfsibiYy3QbtzKAX/XmfrtpTAR5CMJYc073rXCFa
9UINz0ncFMJSACrkIfssLVdwUJvsKVz/z1abBpfkXRJ06AmWFFw89iw8gJCtTzcabD2DtaO8L7d1
p7+UzhjxZDC1BwfBdPzWBPFdV6dc8hgOE3UpMLKpOZ/qSq3aImuEFiU2+echvjgzEk4lBcVMZvrl
Woo4SDRHmXyMYBOZpwgPhkJra8uPhbnpy2BmykhssBzNB1/E+rMBrMoHUVh59S5TgO3hOW8zIoR7
xh1tHfBtX6SLMCwN9FKAooSifVtTS6T4d7c+IKQw2jODzWdZF7wrLfPoiFNw+kr4iMG7qIUSLckc
32oeVoCByCQ8SCNE4TDMy2cc8YhmSNkKcBk+MY80T9EV/6rG53PA0ppbKVTfjv48eqOF1jI8cF1k
MnrSKZ+sJMrlpBH+K087oFBFhMQAkTrSkBK7C7SzUAuH5onF+vcSZejFvU9kVuffmHRP5LN3NlDh
raKtv6xofu2KNFlonLJOAdMsCnY+fjaTHNRtiRMI+0DuWxhmW4DolbCtQhYbWF5xfS9yrk4VCo1h
/AeA+YqME4DhKVm/VQPx4fsw4lbugJg+h9iiXnyZ723zDv7fWpuGPHL9fUb1kH03fQjcolsAtz8G
VBm6Z93mZkQm2qcepE2zuVSAQKteIxBSN2feIOkqY5eDz2xNjGpwKxVZirLycEwRKPHLP+J8/dCE
sk5k5SVrtHsT2XD5kgGe3jLagqJNvbTMoEYP0QwR4WQvF96NNsgLUq2Axro4SUlbNpSuH22xtgM/
KMo2kQC0yJPumK5gerLU7U0iELEihNvYnDS5QMaOpxXDuJ8Nh3NjMMHTlSS1xuUJRtlirgynsEqC
o//ylJJqCV/alR6iBBOL9sfUHlCvBwmV6xuyAN3eQsRfYepO+RntSBYzIfsacvSsXwfVWfb+ZkPC
v4V+gLAozTEqQAgca7a7DVWlq+sJgprsRsw9lL0WkiupoKCsMZ6zrXMJGURNxFXhvT2Qof4G9vez
rRll0J5oE8YYGZpzI83p/AxNafhi6Lad/JYOoAYTQZgzgEEyjJXGGY6/kq8AfbGlux7Ks9H7LfZT
wbqMX42S5UERvfBJfH/ztqx+SsQOxI0ycJ0FA3rQnr3fapamntayZi1wluZF0lSEWuOuLk1qIN9K
GYYSHdVBu72oCaiNN20F/gwIQzi3EOTUEDSKYiU4TgQGRekHZBl+GQyUmFLJAtKmUebXI9Gi16Tq
oBlXGoEaJ7hIz/xdhuubWB5bmvkGntR/vfghO/yrBKVJirTnUZtnTJn7c7SXfBEe6SLnlQIYc6X6
B+n85WsMpmJx34SCyEWeQwgZ4TW1gWi+BG/OpCpcMPr237wWKK+tzgpprS5FYAL91q/YMds8Ob5J
dOSLKztqt1hQEDAtC2CIOMkvcbRlf5VNUcAcfXqDm4DSaxvqMRzAxMPXTUNW9nmwI86Fhrj/jjS5
JQktjuMZ3DBB8G8vnkOLUNkRGMCEMjpHZsxvMC/+Celgwr482lCUSASHD099XgBYVcHoRbeAETR6
JzciiO/8WE7mpCiysELLDSvoP583XngQ6fuT/i558AJlZptsivSLgCs9aQOCWKp3VlN1EkQP12s4
LhRgfRAXfXi+FjO8zZ1ytfszkCMEgSJiyfu9JP4cQRazVu/PXj+uPhU4R0DZdGDrcyLU7eAZtSKY
OnWYbjazwMpJcG5xsJaCCVdS8RFHDI7ayLQ1tBq4Byk54MPB90exCTKk/WZrZBkz0pTgcbmqTlLB
Q7YalzbFMg3HmTcKaW5kvajTDhUMjntV+YgIPYYYfXWoeVtapllCuG07ONditgG34+L9+qkydZ8v
sjfQEVW7qQcxyXKuuEoMVNafc86hQvVi9clUNLONdMTRwq/vIN7AhmJUJjybBIIFi/DlNHmQX+yw
4Y1kK4nJ8uN7AmLs0OecjS1DJigGeD2EC0S+W8RnQJxAmIDX0d/HfSlfvBchesrMVnuAuTuwZdPa
aCvdV+EX/W2Iz6tWGTlZmh1b05hpbcggLgMRjWNobLuC6ssxACzwsNryL/IdfxyUSMKAxN1j1mmI
ZV3t+wsoX4puI9cSbilYF6gXQ14qJKHwBtuu51qPFh3wkGp5hoIPlOTtlaUj+bV+D48iIs1Gdxn4
YaRTAe74h0N5N2oJ2GkaSII7mc0Sys7KFyYCHqdJs1vDkm5I2uCbEg4+5P5C4/HpEMt1CUPMNhMv
FdJ7NeGMPseZWS2E0EQx3gh6YhcUDYyO3/SDS3+9de6R1As9tSxvw3ksBq3Z1s+aF/JW+vyRAjRV
Ok87nN1XhBekFCIDqwLME+AaD/XZMEOLtwH2lO0Np6irNvRfI7O9hkxcrlqWUGVg/UlwpK3NbS50
toBihUbBQkxX8gijREZ/PuYktbh+93OczAOcUVmnc06e2OoJ7PoANHvFfMdMHZ/LeigOjZ3DUTG2
yDkiXlQL/CvybOhYCBr4BL3vNhAhn7T0q/pEyb8v4/YWjOWTyUPhACJifTFNgUbUoC6BnU0wphu7
9FoPFvcelJG5Gj6pMoDNjYPP6NnI9NSN2f/wOmbas+esdCgjIgW1Xb3viKkSx559cZWp/mafKB7Q
LYcnFavDgAGALVm0g60JiBInKUJf1fLP1VO1beE17BMm32HDSM6E4c+A5xip80AK1UuX7WP7Q2eh
p4vT1Slc9EIu5Bh8ACXmEgeUVGsLRkmg2AxkD+sTxKJrwJGC8tp3BdY9db3xxSiWp88rfj7Oq+Mm
H4m7EMrjzSA5PTEv8DX/PFayfEcSX51oTpjXQeCzIRSr3hxLR7/KwPPGySuLjvYGvF8rSTrAgvr0
HYTLE5/AgtLY1qJG2A3egyBoxlpjtZW1qo7cAYjtwAlucS4/mMuEWHSlvv7AWVfjOOOmesuUmBdf
wpCDKR4Ev3AIH6ePuZpNbD2g9wbr0jRuE28yxq+486puAv4Pm4E54gkqvUfwnS+QHI8Ol8iWov1s
B6cQ5dmxZYRFFdpUc0bVJGcI56C4/utzGNIlQ3TKfC14BGToerhiZ5mZdwylyzmQjlZd/221ICqV
49vwiKt7kgDu7eKIcQxCYgXnqJRgwAE2qoSN5hO8kmvw71LlcJlLDsfwASjNI/KyHxaaPyTUFPFZ
xvcbDaxBlV3nXFqCxWfJrIH+n2w/tVtCTLj6R2O2chriob9h2t3X6yI20spvjzIc2Xi6jOosVTTT
S2teu7YiPGqwSNab/+eadmteCQoWRQb2Nh6Ccga6kWM0M9x8+5OP0n/FdyiTIXBpdYdc8eR7YcNl
3vvygaeMBS7TOFSMNdsdkwVqwO8kY+PYq5vYCDUOrHjMWD1UI/7A4vPTfr/lmXyS08UaTHY9jMVd
QLohaNDi3RMRSB5/NAOH6zgfpBellDZia8JpVtPHhDJSr/LtkfMRPLGYXXJzeD6hToZs9CX2WkAM
fBq3dsL3RirNlSMAmV+JjdgfE41Agd/6dqhF1PKXvxCBKMKf6PUCIT4f3kt+r4ZfCuzroeyg3D59
b6XnzJp2Ft1h8GvIR/6Yy6eKOzKdV//U7RykW1Smr2rqMVeHfz9d1q/UYwK3ScoRf9of8mV8vwWb
8Pritut5MNr8Lul6Cw24D/+LH91fV/FAkTyRvlk589wauUw52YAJbrG6YC4x6+dJWWOLCW7t49JZ
8O+FC0i+FXZn3Vhkbv21sAbYhKQcHMzoymR8e1Y06tGbxTCJHmpiih258QHg0xo4ImZwcYgNtB5g
ckH62Dqt/gvQPMuJXidM7O3C4nc6jPaOhmV5qWyAcd2ZWhHqfuOmw38s//8zxJWYsf7+1SGITaBB
4h1lk4/DnCzShaFGxokcz/mrTgoWzOz0mWL2axCXaldvcf7lFPF+YtkQFbZ3OlgSOW8cHfxXoN/3
POxJjvwROGstM4qYOp7ND0KPdtdv4J78wekxy3njgCeNK7IeazgPy7glBxL3pCixM9Mylf93AkZR
slsqlKIi3IzhWOTziIXW54TjO2CLeI23nJFsY4BVUaG53TubsjxHeSwzv2MGyfWSfIAAfbbSUydw
TE/ACj1LqRYCZ74BTj0L4QKBGxdSa4eW78vtli5jClYAT6yhHDQjXrd4zcI7uQjsPJ5we6uAbeJ4
JJNTDpqyss9dP+36W2FBiHzC5Ey/wm16tL+xA5XFYt9yPdHPDKDKaaogSUDLI8GEc/gE55M4yadt
1j+4DkVb8kZFy5FyMLq6FMnoUdb8pY9RSkr1LLNPixaUxYAq/oBCs6m9SQBZXuR+/G+oBl8oWZP1
yk7fxpjeGmZJ/dzB6QQa53B1VF8l8VkXrG2UcsidqPhE7RGD3hW7q64N5q0POl2ZYIjHFF/UcUan
WsKUuSlXnNuyWZBthvW+5/q1ZApeDc8sbFOTEhfSvL4OCpq2Vzpx/1PRTpjS6sNGNh/Jpy+10ahP
YUVPruEvSJABt7DpX97wuDsJ13k8nvXAc/34CmuYOzZxI/pf5VYsgVb0lk/S2SoM+mHaELdb+1Wl
UbFJ3HoXXc3wzdLVrYGfDO8DPijkQ2mUckw8M2EboM4jAeJ/ruRhngyubKobey1A3YH2EAlfhRsJ
lbAnjPfWozNsBLJpIC0eN8zFso5A/vjueUFMCerPt4PF7l5uFO2kimphGjCm+ng6t2Y92sTZqoaf
CuBwp5/Sb9RmuM8GlD98Qho2UrAi92PkhfGfji+HqreslWPxhqHNuBGMBoaJuUmNcTpcWws5zaIb
U89nLcIQhAF0Jc0ZKf0bmevSrS93CpqtsgPP77d1sxLxM49KYUXro5AzqBO/Vg0a8z1Dw+YtiN/a
6YGM1UN8mpoT+foe/7ZSOax8AWmwESsnSFcUYhy3IVsgJYaXKaHrX1ePbD2MfRSTOaAf+oIyHiab
9CPONnXpkcJRlYitUeLIamP1MUp6WdixHxVfJrncUH+dYFKR0gigUm3dm/Ng1NqDGcYqjq2hOCJA
bYDfQhRGRDcqbQyWWhbu3Ukshyw5lhffcxys8+xC6O1X7/smN+S3ks2wVJ3wjaCEg54HbOW6NqcK
ujJUTGRXu878fznDzEeM7XCYAV3WhszsrjQe6jwXPOg1fLlAVHITViOFpmKYg2Vl7L4X/J6XFGCg
/SqjNFzJRjRcMEJ+anEEu1DhVcl5oFXrKJ62jSrQM2JRbrZvKBEed5C70N5adQrNzy5+LZIDF+ly
atPvXzCHPRwEPUCMp4bXOKY9boJ2Xru1cxpdW7SNa0lEvUWqliN9r8HS/eS1c2LDbcrq3JnH27CK
yJ0rcT/4rO6zUS9rKcAUH8UVYEZGLRpGMe2pMpvgvSAVeF0AAdoTI4fQjNwl7kDySUr9J5wDGv6K
z1xVnrGdVUMkWBzTPaYbnD4CS+f0b37i9snTnxFTPEO4DzGgMouuscrOw3YGyNZesR5jYwCMo7J7
9mGFcRnHjh6chXLzs+rKrUq6pOWDG8BwIPrdE6CkC69q0OF568Ctgc0xe46mQZvB9rFaTdvj3dXs
AqjV/rmr2u3sXmdu14hgf9WaNCQ3w6W6HP384Oo+ZBjzDT7oCFjZlt5Td9eS4Uw5wUYavGtrvFx/
NgoNeCxYGWGlVKGQ7qPGsuJQWpQ/816fs9UKL6j2FNusElypuLvIbjZDUo6zME4DtKgWzJKAIvUA
iTJgUNq/eqM2cC/hNsaKbK3oPvLsygfvdfd6E6UdtocaT5HwowJn6zGvzvRseezzm+O2MV7BAGPj
4HRv0Fgxh/UvL6+tqj1HpEAHJYtLL/hogD/Jjog5/k06ftO+tGca4EQhR894OqRffocFyH8sSHKz
tbl2SZ1J9245HO384Y2/mOikIiV2b8pkO8ffGsMvao8apSeh6nYjc1V18RnKjS8UKm35lc4of91b
zY7voWaE2dSij1Hzu3rI3LpEm/mDQ6SoWiOkIBcFd7v7f2l8dxMrDmM/NAaLqhtPR8C+Q4GBSsVs
9XmZ6ZgHzkHWJYZDz6ZQTmJoQwR4nDNV2CqT5+vfHvezJiPON4cD1YNyDcBD0CC1ehA7Fmg0JAJE
uK+6RSVHlD3/rAX8JMl7axbYA6e0Hf8QbSrG2JET05y3cKwHfB4fL6olEigxusqFbpXInHwlhNON
XK7I6NBn8tZyQ8yq9fVfgFHa0w1ncNWDuRi43qQZfCl7Slu6ER0tc97B+41Pkg1u3EVxIyzgzVyK
IA9aSJJm6q+KjR9imQA5bb3AXgOpDarFkM6TEK50AY+RSYCeUWTpXw3uzZ5jUwQdi+0mN3BVK0sj
MOxRU3VPTjJQ83gY+QhUiYSlT2sFgngYUseu8vm4V/H0fijbWUJOV+0/PG4UC3F0PJs8WtvyVs3r
7b50QK8Ppc3o+8Er7Oi3PHsArw8gZmiK8v5vaUWcfDGtkOYyf42Z8p+u2zvULNv8DLttGAxuVHwj
fE/SqTYBtw+XuivdWDcKuvOAq6PBLl3kKzEpLzjokrWX9UmMAcTMtYVz/q6QlAx7lVAYh/aGFJiM
UiGDxIx5aY1S7LDzQdA55qoaJwvOqJMqqE/wViGzfn9fp9v9p+lLtkWjdGsDNEJRo5m5U1XGMtQq
Uavy1iPoM9e/6XnOhRijhyectwl7o27RtYLALjoqfxN7Wp0Pi6bY8bo+1rQ1/QH55yhgNFU1izqt
y2V3uUOnmiCKMXfPvky64A39jI+1aiJI9Ue3cg7a3pgiVaaEOAEnXUA0AMEpIqBcabYTZdOLACNc
o75k9jINc47i6xjzM7W/y5V9N1/bQkbziuhGBR2GIW6fv24XLPGDWAYM4vWGFpw4sc4gMWIP0Sg/
Pc7XZ1W/5Q3HT3nC/gf8AK/dtdeRAoCYzgUggFL+1Fn+E4VcQ8ipssNGD/CpgQUH38EW6KoXKcHR
HI2TQA7s6jbzMMqKMFsWvpvMORynLirn56+t1hEo6gkAzXj9at9UB1Tk7SFIhqncqWzGTjq/JYMB
vB6ECDq7uFoyju4UHXSNq+KF++qFjUI9JrjW+6AKh3qW9/mtTinOdSZhNOE7hkN5tdaZNFoMDKwI
OnolgbnqUErNZuoTLKFbyEwFdY7BOfQgOX1DdWvu8M69N2ivy7gztLS8eN65S3GOVnx6rUZkRMbq
WByYdv1w3G6onfIR1wkpMamuMSZQC4ZePCcLUX4bBAQ7zhFISPdrrAC6Guf4mPRWek7y1RzBJxvf
Zm7gX42hISRLG64BbrpGCNdFwQqeVaP+SnkhXdJH6KpYXbEIWTydrEa6kk2COvpqvdruP1I3ptua
Ng+EnMsa2h2gw54QvHqdZLiT6n8mWmM4u6Ooac8ChIUkAZF7Cu4hlGJY8Dmz0RTay8NMspmRIChw
raMwLwGndN9Pa97PElARW++Jb2gUi2S0D1YBWODwYSPODU80gJH6/4h/AnppoyGSp/C54h/DR5Dj
B2PXQZQWGc0Rb4QqQrTQbH1FgdBxqanKNEALjfNcUgkGTpMtkXQZ6f2fslyLO+5Ro+dopKLfH/Is
H/HvUGUtaw5phgDRtopDfxZbDkm44KagFSI6Yv4GMlJ6t2E3peRi6U2lwc0zVveLUMZkw+N7jixh
nE5AAOeXlA+kMJPpYblzh7i8TqRRiFLdwGjyD+DE62o16van29QcnJIpZbpgCYTt7DRiBtOWMMze
zR/i5cpEseYFPfpURnxVLKKVMAPoWoellcLuA5H9u9wck04DIMLdQF7ErtyLToS3oObvtmZht4RQ
xnwHZp68RxKLPCvGHXJhjeaCR0Qqe6F6YZB4D9o+/rUjDUpEbInjGsSAz9VObd9TEDiV1bvx1I+C
4rCxsK1sFLqPkEIYrpKafZgFmY4GPTyQo/1kH7+0ct9fCmFbwSUhrpSBcu72iRI+ctsNxevU9oJD
YfWRFC0xFGqZ6Pc0Gp9zjwLn5+dCh3thgaf3hUq36pjLhdeyf67Z9gMC9Ifxi+BMKebO0nnXzrLb
ShI9VqVZStiKZHR4HcL5KvNnLGcleMOBr/XL9URS5c9ZfA7eIOFuz6G10jABrQIq9r4VjmRdiqdi
x9AhLho9r/m1CVe4GKSIxSraMzZb6Vky5K7l7qM9stxFltdWf7nybRAAql5ZMLVTbZzk3PUd6IPi
wsdXjFMTt47uhE0PAWB2uyhMZl0cSue/7BiCwXXavAyuaBI1TNjpU5g+fpi56i/f91tdNJOqxZ6W
WdXUTM8O0q2xubCqe5TWntGDL5iBmchQx0dbUOLvsAm7HPj3o4aw/daBjGCk2UzB992hH/Km5QpO
zT4YLl2sFqRQOX3Bk7Nop/bVsjSjLpZyJo0wd9Iwr4Vnn4skY8WhIxrSGY+0e2y/vhemKH4UG0P9
r4QFJe8wIgXwbw8a57LIUvzeVg9LhcwFs4/PNWJhBKefioPv0ucTtWvQdk0VaD6BjJVpmdIsGuyy
S5A6VZS+C5SdW62t1/ado6YDOtSvo4O/1Bv3AIAC2y+HqfuSyjJE9c3QyApDLBdb+TWGpGGmoH0K
dDViM5hv+EXXU6lzamZTPJhRujnkkAGPBOex3+rGA24nwGyU3pFM64OW+Plj1oyWI60rQtolpjFS
Sk2dGM382WDaoFLI1ihjXYEysNNIdSjtO3RMVxPnBXubPALS0U05A4ls8hvsXA02PZQRzuecn/Pk
pzpnrlKXMT1mzuLqdu2VU9hviT8NiPm+/6GUU7SVxTC8W7dZAcIspJnomJ6970GdxyBHJ/1C5W8R
JlLMyw5Ogd89g7wAf0PbKoMJg9irycNON7FQ9jUp+VXCq0vohPZybI8C4XR/6sraUnFcYi5PQObn
50Fy9+5A5I3uDJkdFb8MxxQYobU3sf94m8gm/BroCPMqfK4eO1fk2KdBjJLoc1V/qksjeam9Xz6A
WFK+9BeH7t2Fn/Com049cqSmoUxQISqWMmb9Z+BOrnOQu06E0OOgTt7E0cU3ioOPmfg4c3NLZklx
jy/lFbY0pi9kSE9gfPVjITp7eogBf2VhFcqxWaihKMyRBYZl0hjO1cCUg2qqvTVezLn2S3sL84GZ
Jk/joWk6IyeGItdI1l4BTR0OMVwCPRbOKn5nwuE9EK3eDHSlez4xIn368uiW5dQ5kOeF3VaWOFuT
yVM7V2qigAOT8vN0dIqrlcxd8akwY2YRLEMhOaVaRzvJFePsRuNJxaiGin1/MCrAHsXYZ0PK+hRy
thLTtSOvZyDU0p9KnQPeYRq5jFpbTh9V5+q1mX7+4v5ZpxYZgeUuLvC7b5o5WATxG7inS1uh5BH2
sBb1YWCQAVJpr4IIB6GRmVLX+EViNSS0CQlQ+GNSipnXHiYcpTMOw03v0vNteq62vWA+c5rPgybW
E7aqEw6VnqJCOB2RAEPgQwd0CdL3ahOreZyPa5XFu0Aan5pE2/AzHycPM7Hz9Bo/3xdHL0xu5KeT
QY40h31A8j/dbWzTT9Nm5K9WftdpqRwOa5/FLsyrgjnIsXP1EIkcty0TmL8258AVttClNjSkBohp
Dfrfdam0OI7wmTCd9UWpJ7jwxFZEozHblwrrXeh2sUXBG1xl5vt7SpNdWQyzTrlTm+1GmPUK4K3K
B5l1onjTOcsbBulca6hUAlzRtFZ11JES7Tg+usQ1Q/7RmUwO8i7asNt0BFycUl8GMMm7iXIC5DSO
EveDAIeme+vv/gozRXTqm1Aio5IrdnEfQfTLNqnBMLAQioqWWh7Bu+UMQmrjIuUzJPIRoFov/Txu
fbmyHrGUdzCzNHP1lM8tKvU9ZV/tiE6tkrEUvVNVsDSM+cD1hKgmhxIYuzW9ArDWnH7Ys6q5VBua
sjiPBmX0jGqC+mcLumRNh8L1HjGOX5WArTtGk30Biw5l6PM2Uj+RbWZNiEj+OtxHZLehFDRRIkSU
wxKpfkmknug6ABrDesAbAT6Wyizx+ng/sBd3gbG2gIQtMHrKRbaZCwEvrvbmaW/AMbAusIJ8IgTn
adysgZX4/8dlG23qU6jSPTT4a4OGFVjPwzXxBGp3kbBzNgFgFZ2OlJRr4zYric8kxUrvysapiVAx
29Qa9zyyOl/aihj96ws/zvsCidfv9EiXEBljXPv3gG/myEyuPO+aB870kgPWHFg5RIFxBRUd8DNh
4pmHz97cjuQUgXWDbfJ5GEbnXbBSHgLTRLcUxqoycJAHSCNUyLRCxPYokvsEOGjHZFHo9WlstQIL
mZSkXNTlvN+um4JFRhrOfm0haC2EoaiBY51C5KzRU1yWgaspLM8Mn5YRES1x2+By/3Oo2RntRNTO
Xm7byjvCe6uN/aGL3o4VrBjShU4qbCZ/IdRYOrtB646SZch/K8QNesKWmpS6AZp2SH7GxH8Za9sm
mU03E0pfaBKIrQbrlK/f8NfWbvEmrKqX8sQISfAEL18VFWmjZp1xBnwkyUGhdp57Jh27wI626c7h
IS+pm9BzWY2KleJEF8LLGwpfwOGTEMnr2rxXdFLs+RttiIvFFgv9M/006rAOdvrgLnKE0DQaZkNV
NLGr0rS0G4WYSy+aHWBP/2sBGDwrw1TiBBaf078t4zjeYSp+Kfor2kwtfsN+frr2+ZnhQ8PATWUQ
xxArw4nMAPPCbxelTlpw9m86+Sjgqc1njET3E3cxxaqCN6YAwpFGVHCOmnxflEF/Ppq8gFEQj3yB
EXCnBpnuLaTk611c+wD+MFeSEXeeHQ5+yyMwSXqsvnBi5WLq1rXDgIaW7dz7CjkSq4jP1ygKWmo3
CfmgPxOrRTEwNCgelEMJLRiMj70bnRmTXf1+ai+HyUMuTiaC3lYPeqIaN2OROyCouTSz4d7Llw3F
+/G7L5hutePGNH6Zu4MWBe4ENQzsAksNGe75rHDFbrzXOeF3DI9kxGCe00nmbkt0U+ppUaedMWJH
x0cqL6y+pegV5C2147EUzuXwuOrP7je7p4vFPNJ3Ns9paTneQnX2RRFkzNhzYPthKSBLjCJuX2uY
r+qpndiF/mdm/Ta/mhpbeWCAUPs6/qncnX1V0ltud0OOeoRTLo0bSmntGOUMLBaCm/XRCAG9nrqA
dgCj7Sk3qTf5GFX9zD6Z5DEeurdm+nSP9H7O1TDrGc7ZXOA/DsA2kHq47TQluEur6As/vCc/eaDq
+okT3Wbr7GNCHIveauiCpr73AC7CXYH54UJNWXcv41Cqse0ldE43cioGJnho8QKIcDxdqovCQR/y
RbYYnPIm1m3RfypeEuJQ3qgJ3tEGfozpVbVj8aYyAd3z44Bkb31PgKLsk6BX32S6WGie7rvS6E1+
R7D43S96ovH5S2a3JPelWzbOvKVu9x2LAAbMvFnZnYEmdNTYd10PPOk0tcQdOkF+kROt1YR79Uff
7LwXXOCWqTbv6IhksQYsO2ws6q2d9/1+M7moKwL2Muh9KyTNfFu4q/yebzAP1j64W2FACIYO4WNF
uVk7FoeMD7lGz/+HrwEK2h33ap98xJdkKHq+6QLa9Ea+7ki7R0wsNs9zn3iSMQhMIsh/Y7VHuq97
Zi0k5vR4uWIu85yEDfs04jeez+piUWtsToKgp2h8hpmahk67PohSPLlYfdv7kzNTFuThDqcYJg50
uSeUn7nu/IZTu4EMmWZjCcQoo0v5imoGBZfWLsaJUxqYFtaqQqFV5YmQecrn+XTdajIv/bW5wweT
YWFYCgZRlkWwj+u+oe+Ey/HdQUsSlxyzCpQK4FTe9IoBzL10Gel4mnvWKyxcmWUhbmMn9NUYEjfb
JYL68eVDJe9aO4upnWD4ZPvlEwCxzrKrX2zRqunq81AM+De1m2Dlyd88+5jhmCvWS+2maJVJMuPu
fKGWVxNIM+CM6lx8usLC+hmrt8Q//F1B8G5uYE9wZxRItwCoGqqkNzr1LtZL56uejDPAHHSrOdza
9o+bqpf/VnXlEn9a2L08hc3NH2GoV2ZHlaRCh5I3MVU95eah8X2d7dKGlOEbDCojez6qzYR4Hoqi
A0e8usGr5w4883xBqywIlEFfMuOrMJLJU5kkQAJdb421rd6P5RbnqRkivsjT9JD6dp+duLjUFUFQ
ndG7O+NvaWlYR0OEacCxW1+WKI3SZfO32zGTx3zm0inoQL9nm0GwDddkDokZ6WVG1IhHPYWOGpmW
tueubxclMRD9EICnS2e13Zc446diBiIsd002R2Vxl6JXyKh7VRkyp9y8VDNOVPniBwwI3HU8YKp/
Y8pXLRGYrlrsRI6XMhKX3AvHzvZMnjwwUpCcEB5GqeEIRlLiLZ7+ZpiOex0mLVM2K6e69Gf/yt9R
cV8N0ERcbWDNojYzU/7Rm131J5W6gOCQwvejyTr2Aa7XHL+r7T+DcJniAa65wWC3Z2P4U8uw3Rtq
FeiON2Q8v8cUuhFComWSye5R1tcxOXahW5v2AYNNcNPHT6Z4Loe/VCqvHETFfAcdQLuH9qelsUlQ
yjcrcBJPOetmehBdl81i/miJp74Y8rawJIW8uIGnZhOSniC72gxMFGgAcyUsCmF8kn/bdxRkHTSl
RB2hFZ3v2mZJLclOyJdUdyM+rqyRCOiSROSyN3arULFxGKNU4uPx+jupPTXlgqeI1L+9cKeTm2pJ
GoLj5DWLYi65Vro2vQxGVdEbwvO7CEq5vvbaRB6yIcd8bUpyZtyAwqadiYH4vydmWaIL73sS72+X
pPsn1sQPskZr07XIixtKhN5jDSRbfE9w2jWs7fRKygXuOyPrQgP3bP5ea7FOlkWya+a1OVRVk1Eg
28rDQv7i+nRLLF4T5SfIeavI6sf71pAR8wUy7oAf7JMZ0k2jGKsthD2KTPA7M4gF57UEAmPGaw9P
mhZa6XLDnALsEGeCLgB6rINL9y/hDp3oou3F8paFpjGLAtTQhnYMyLA/bz/CO+vK4/LAMIZhHrYp
PhKq1lbC9jFxsXcwZDmsZoVuxOv/FgsFnRn5cyCnd5U4wyG8xHyfv+Tb3pkL1uTpDYYG9+WoCKXU
dhVPB6SNQbUt4UmLUNuTkLLoVOgfNKJHXibyO9xMpBAKbOrHQ4cweIobk/rGg6Yedm7LuJdp5a68
1eMS+8W9ziPWUTLe7JhV0X8B3+nXZJyLZD9mwPXA0RZHm57Cq4GhsT0huyURb/PYCEOcWzsg0r8l
HKOaz/oFiofktCNM6ZET0EUkFJbgrXVjDbNwOMsVI5PNEdF95rR2byqXgE355BxCrfTTHbBkDkxN
5K477cB1wpO5SQPXgjQgDeOQc0BtcuAGJRTMXQ/OTsbK+b2w9P7dgiOKpzji5vQ/gfb/YmGti/yw
D3v4DyhaDc80CyMqhNSIvxZg3wr6zu2mD1EdRtymHLg3pObHErTisFFCNz8OVAtOgQsVwdQTQtdO
kaBMdhgcxtoSLsKU3hh7ZON1sNdkSoBsL0VJiv0qFFNMkRja8/ZbzOOVVBd7fuBHVfHg064cD4qB
j1yBudtHIh84R5tuucWINFIMjZD4gxAcue2IvTkw4qwmsjjMrSsUeZuDzI1VBWsMT13U/Tv43Wod
yHsxw0kLwOBnj4DDLdUOEarYx3LueOgJCMj3GcfuhnhFMEnIKF5MLRHaqOmcGikCTCZ4ElKPPoMd
FfT7rgibgzrUceFod0KfH59C5P1bRzGFw9MHg5qpVX4iYQ0vIy4R9IqWhYpyZEGwiIw9lc4016rq
TRWUj3QoOx9p14IMnxMOlpzFKk4sH9EZ2tk3fhYTJ9Rct9m8WB7KB7Qaex1hAJ9PjyYBXGBRBryw
mlObcT9JmvAoMyP7dIeotVGv4wLsoPTlDg7wS1reAceR+jBaG2ux21u4X5KR7Hy573VtFdX17HLU
+TTb8v110OFTJal4MUzW4gr1OglBRHzO3iV+1BpUAJyo1BY/8Ifkbz68o5yuozNeNZCXyTibj+U9
em9ut/P7V98/BGeggSY7LIZK3MnTxqruS2uwQWp0E/Zsj63lmjTSL5T8zuvEOMGScFnVk/0BRzoT
WSWWGrURVIXuEQIEBxaRRXVfR3eR0jsSNgwl2Z9mCWKdvwzOQm9MTpLSMICEoGqlM59JpIDZEId/
Y9Sq74YH7zr63l3mTYybMVVORMJu63ER1W8/4K4sgdQf5fuuRuqLceyh4IgVYTPfvrNFu5J0I3eg
Uqm3WGdR0KzNyZW50H2h8Zd8Sr5dBgbeu2WnEwGEoqNCtoXuR6mJDikni06eekj+KX0aIH/dARiC
qnaDs/beQnsMSXarTR+XVA8eQM0buBLyqufZbNfd3e97WSWA29wXLCE1fsTBMq0Tlp5Jr1rRn0QS
v58xLaM0APIxL5hCJoZkX4ENgot6W9ueDI0kwxN371PlK0CPs85FIghg620JlNJx1BPkJQ7YJYEs
KKSffWyaSxSEWBJxmc0g+RcB5a4X/qd5noIW3qk/mERT3DH9UL36uoafWxl2MWYyLUS2mmhvHErv
dDeAQm3yNgGS/dBekCMJ3m0uJE8EUOKA9EGipkx9XzjZJvSlMeGcCBMVD6Z/zVJ9V7lWPrgBZLF6
cveTmMeYNvzZpg84ByiK0iVuBQicN6mhTjNLm7G5qCbWgM87qsQESF6J/6xsRaIyyBvMCwJs5OiZ
Wo1MAAELxd5sXc3HeXR1Mmdik5p+aAkH87Eob9iJyFXwkF8m03abX4HuhJ3qhh9eaoVSBFKGL+53
pVVOvf6GVnG5mScoyqoYVk5R9R7oH1PE/0WhBCy4QUw0tFikI1bgBB4I0N9fGq57WYEH3wQhg+D8
SmzGvF52dzqKNwt1k9O+ePKIuL00uJ3VU/oA8CUQ4+T2yl3/q5kcOCISnJRkIxB3+1Hxu2yVwag8
Vmmzid8N20+wyMLcMSlexPGFOvBx8dlHXWI9HQ/ta6IDBZkJ7vEKjx5W7DbnsIJf3A5sO1X6qaPX
ZBxHQiteKy7OpFANjC9E2sHEAT5h0T57SVgIgzU3jqlbHq/6uM4YQjniQVoo1i7zXGzD5WQsZqdC
zBtrBrmiPzk8Uu8jnE/2OBu9NmD/PdrP41gBt5FWREUzZ/4mMCLVeWT1qq9Cf7NV9q/03Y4CdsIw
dRBgnV2hEBsQKgsTeb7F8EWBugc05AlBBj99E6H57zAtNdw6wnqvQaIMfvjlWc/Czme5EKXiBuW7
rY3QY2+uy5JLv9e2jmwd3RLFNX6HF9i3bzpNXwgKAtd6Tq8UY7Ed1IeT0y60NHtNv7GZyTPFnfQD
E3keo1nUqsoP0ZuIrV7C1d4XApGGjvzIYz5bzDucrvKHAXLzD2t6y8y7bxagvu6DLWCqEtTuuWka
cOwxv+p+NOP3QYOb/CBoRU3kNGklYLZqI42KGVpV4RyJIx6UFveApL+QqAoeSGwEsY2tKdOAcWN1
h8hMDTM4tWU7mvEf54oV5KpY8P0cQyeEXDFFdETD+J+wOIIlOORHt29UblZu2cas5iemUCLd4nvs
1jSfgZfLYd9AF1/WyJJw2yFwnTUZiGKHSM+5ieMyNBUb/P1A874+uNksJ3hqowDl8zXYaxIPK2gf
YqghNd9+DYgyxX6dvX30kQ8NnBw3vQ5gCGsjOJGRp/XyCZFkTLwdxzgB6W6F+YlltL+SEc/F+Gf/
9KT9jixpBrCwNm5+/p46pzlX3xSHbUY6+wdc9f8fNwy+p6nyxIbVBvnFR02Jy4dduVoYgNLE/FHx
BPqEcYe1tq8Q5o3AoJ3xrVvWTh1gTuME6y2EJb/p9x8tCNs+8gEldV+Iy5/pHJPukthK/rN6cPco
yU7MvBNTq0DW1W0wkJuV3MvqYWVaUD70OVbWp500gYWw5yA9ofVvxRw5XCmVVu09L8EkaywnOIN4
Q4cMdGbWxXeWor4ZNW5NDwtslwRoybeuVw0LLc5BxRO3sOUG8k8m/g0yM0ibF54pxXwnf1ags8Yt
aZGpjUDqNtauSoHbBBQY5dtJLKFG1oaKGpZwVS+xNavI2EeflfAbJDq41jl0Mn0bgyqWBSwrjlnR
kZ8xBWd6ompskpDMKam9EtEjzLot31Q0U0U0/CqosFawnpZpFqDDCdNS7lsqK1K4p1CUZ/uxCAr7
G9hIHOz7M4tayRERbAaUQ909OHAPlb8WdOQvzouFuwASgncGDIiIo/t+cqB55e9R3kvdirWDzbB8
inFTLlX1ldj9O3xjzZGy6x9h31iP6v697JglaeLyYEhMgYo8Ou5UY9L9YdltOn63RZ6Ms5sFmUZE
Gs9ZC1nNjf+hOfTOLK8gWsW3rsghMO4Y1nrFx848MyBXpcLgr5Z5tHknHmHcgi7kkG0UzO7xzTCM
LhqyvilM38o6BAsLFByKNjpbiQlx8iLIsgK98lc6mTcfOCCoaI3uR1GqbfUZmpGNY/CR270KFcNG
LqQl2xPVyt0Lp9y7ZJArDOyBLYYpzjQfviNuyjEFolxBPeoxu4HPCgqJggXfVASUlGGbQuNFIfMM
8f6PQaItIDpB79NFwGy6AD+PP6mhxuDscb5LSgaj2g1JMXULC98JHhqGGfq/qPwIw7wWxj0K3j+t
vTSmDNRwGy3bCJec5QsIRxG0WZI97rjWJdocmmdMtlaMnZ9R/PKHl2PauWTnf+AFGYbA4g8ri2uQ
MAEQnMJjpmHk83wBd3Vjz+Qd5QEJakaAxuepyjTjEddgZlqYrBHehYCLkUOP8WruDn2rvDd6DSB9
syFZdk1MFpUjWZUZ+1+l1NIigQjclz3RGbOJYLOy8zRVkD1P3QBh1bT8+x2UpLI/7xXLXgmhqrQC
5NIz3ruvacNrHzxQr8Kf62KGJacmk7QymV5zCDz9qyUR31JgCgdvmIVRuvZYNxiW5BTP+NztTLsN
c8Rlfw4Hw6xm3HBc8RZ9XcbXlNHS24k7VoNlb6iztNcGaXP2jquYyaUjuV+0b4jaWveptWuE19+m
tVm3PqFpI+IcRNsUxl2EsdNP3feBe+Jodrstxo6v027oyGA82hADONzF0l11nR8B2q668zshwMfu
xYctVXCfQ0Nn9nx/YiP8cgLt157NgZlTBSBPLT9diFdwSVLWik2Ah4qnCKA9xA+CBM0THDcSArYK
RzumLyBhUDYaSw6F8+JKg/wIMXG5b2D6UZX1AT+y/4hB8lJmu+aUXPBbuZs7AdkdeyR0XeaEimyz
wjRk/V+Gh+C/Kp8FfCI/95c3QU/buO7OMFLPBefL1/dZ9iHgeRqEIIzVufVbbjgQ8YS1nSicvpda
z9eK80lFaTSpYTy7yQzpwcS/fnTHwWBFeYLtGtZQosXAim7F80dl8hFk5ctuEruvP6GIYOh8QMXK
fh3Cyp3M+O2ST8I0Kn1c+jdcXCT0d6YAfwdZfIQu9zrbl3u12OklCZ1Xn9Bb3WpiE5weYW5xgxv7
HvlGe9YrwYE7hJtaYKUTLv+SSHbO0i/yZy5FkfB5Lkhpp0ilSL4rV8CHqN2d0TZIGZebBQb7sAv3
MTZzl5qseiOV1GV5emK9uVEF2RECPJjHJ5UuzDqiq7/WrFm8pjaap+23W35acv3+8OAzJ89hhaIV
ELqIDN2OGnejsTD8G60uv0+31j5K/c0LkLcwzlcN4TUR0VS/leOTkV90B/mFX3UOTlR48Sk5Jy5P
yYXqrqpKwSvgbl0MP0FeP1wJJHvXwJkx7FGidgm4mBzJ270j4wT2/tHzL/6p/6oaTwOmeIKkIb+R
7R5yuZjez09DulfBUIwSFMHj1J7hKqqPML27UucihELhnBX3cz4sEt7BTmP87JtGLTZWys3qF0DS
Ycsqarpf117mOqiYeKoJWVws/L7ve6YmS22usVV9ie6wS90OocI0hHssmmXeRllr2Ks15yKlvsJ1
fPVSFOeUmoM1ACW1cT6lZKQ/HSN9odBJ04UhdT8wCa+IC8ej4w5n6oT97gb3I3TC4sn4Z83PqVgW
jcpkXJqTzA+70UonXEziUeJ1HMi0k/kDFa9aSxo98EnIt+j6g3EgdGByjz/754Z7VbFPpQE+8F8U
jsyG3s2Hl7Ws+Bz7AfgrLnJYuEmeeeFaJZnYCJ4j8x9CLfNDoV1pZGjlaXdA6JNVd34AAF0U2+/Q
kYlqAM1CyDzBEJ3+/h4ESvGFRyoH74KRCjmoSfIvVk1KNZubaVzVJDFY9/YQZJugWegalRuz9o0F
zcdWYDcHL8DzuSHOe6Yv1IYcZyrUj2YCkqr9Oy338dFrzFopEJs05fz0CMl5e5OLAuLa0RlT+erY
T4KTqkNNdUpwdvqCDJqi8cW685zFYGhZMgDQPmFxkgsDjadZo7odkVeRB5EJA0xIOoHUqYJv47sI
WPBKZwmCJLmxX8Y9K+1uZ3TGIP40JtKRx3U59w7BiBa7jeG7choR/qzdFaS/Di5MwhPlTNsHEhok
etQ0xRM7LETygzzXTb4Rxw1UTpzYOJd8aB3MECHhtPq1t6B8a6vDaIFNXhAlsDF7+PFArdMkTQBm
KJyuagdl7C5UcmOZdA+N6Z826IlR7w5Wj3qL8PfHFGm6aNNVEgi/LQVBv4HVVBQ6yCkdi1uhwvIi
N33cao3s3nE+UB/On4SateyxtxEhRbLv33/MZVxIJr5aNwUyrauuGoRvTHCZY0BPlhklH7GPPBR8
fX9fF5vE2XfDRwL99z6KhC9ws7z8vqOHeGhDhuKJ3LsiAXP3Ci61C4sAwtNk+BcGe8n/ocMJxbAF
z41jBcVn18nRMHameAnYkdBtG0CtxnYcOg==
`protect end_protected
